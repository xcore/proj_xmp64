*
G04 Mass Parameters ***
*
G04 Image ***
*
%INV:\DEV\A005\CAD\XMP-64A_1-1_9.CKT*%
%ICAS*%
%MOIN*%
%IPPOS*%
%ASAXBY*%
G74*%FSLAN2X34Y34*%
*
G04 Aperture Definitions ***
*
%AMTHERMAL90*
1,1,0.0866,0,0,*
1,0,0.0630,0,0,*
21,0,0.0867,0.0197,0,0,45.0*
21,0,0.0867,0.0197,0,0,135.0*%
%AMTHERMAL94*
1,1,0.0628,0,0,*
1,0,0.0472,0,0,*
21,0,0.0629,0.0079,0,0,45.0*
21,0,0.0629,0.0079,0,0,135.0*%
%AMTHERMAL96*
1,1,0.0943,0,0,*
1,0,0.0708,0,0,*
21,0,0.0944,0.0197,0,0,225.0*
21,0,0.0944,0.0197,0,0,315.0*%
%AMTHERMAL98*
1,1,0.0943,0,0,*
1,0,0.0708,0,0,*
21,0,0.0944,0.0197,0,0,45.0*
21,0,0.0944,0.0197,0,0,135.0*%
%AMTHERMAL107*
1,1,0.0943,0,0,*
1,0,0.0708,0,0,*
21,0,0.0944,0.0197,0,0,315.0*
21,0,0.0944,0.0197,0,0,45.0*%
%AMTHERMAL109*
1,1,0.0943,0,0,*
1,0,0.0708,0,0,*
21,0,0.0944,0.0197,0,0,135.0*
21,0,0.0944,0.0197,0,0,225.0*%
%AMTHERMAL118*
1,1,0.0786,0,0,*
1,0,0.0630,0,0,*
21,0,0.0787,0.0079,0,0,45.0*
21,0,0.0787,0.0079,0,0,135.0*%
%AMTHERMAL120*
1,1,0.1023,0,0,*
1,0,0.0787,0,0,*
21,0,0.1024,0.0197,0,0,225.0*
21,0,0.1024,0.0197,0,0,315.0*%
%AMTHERMAL123*
1,1,0.0921,0,0,*
1,0,0.0686,0,0,*
21,0,0.0922,0.0197,0,0,225.0*
21,0,0.0922,0.0197,0,0,315.0*%
%AMTHERMAL135*
1,1,0.0708,0,0,*
1,0,0.0552,0,0,*
21,0,0.0709,0.0079,0,0,45.0*
21,0,0.0709,0.0079,0,0,135.0*%
%AMTHERMAL139*
1,1,0.0786,0,0,*
1,0,0.0630,0,0,*
21,0,0.0787,0.0079,0,0,135.0*
21,0,0.0787,0.0079,0,0,225.0*%
%ADD10C,0.0787*%
%ADD11C,0.0630*%
%ADD12C,0.0550*%
%ADD13C,0.0709*%
%ADD14R,0.0709X0.0709*%
%ADD15C,0.0591*%
%ADD16C,0.0866*%
%ADD17C,0.1378*%
%ADD18R,0.0394X0.0551*%
%ADD19C,0.2756*%
%ADD20O,0.1575X0.0787*%
%ADD21O,0.0787X0.1575*%
%ADD22O,0.0787X0.1772*%
%ADD23C,0.0315*%
%ADD24C,0.0157*%
%ADD25C,0.0177*%
%ADD26C,0.1181*%
%ADD27C,0.0750*%
%ADD28R,0.0750X0.0750*%
%ADD29C,0.0079*%
%ADD30C,0.0157*%
%ADD31C,0.0030*%
%ADD32C,0.0157*%
%ADD33C,0.0157*%
%ADD34C,0.0098*%
%ADD35R,0.0236X0.0236*%
%ADD36R,0.0571X0.0453*%
%ADD37R,0.0453X0.0571*%
%ADD38R,0.0394X0.0276*%
%ADD39R,0.0276X0.0394*%
%ADD40R,0.1280X0.0650*%
%ADD41R,0.0551X0.0472*%
%ADD42R,0.0650X0.1280*%
%ADD43R,0.0965X0.0925*%
%ADD44R,0.0472X0.0709*%
%ADD45R,0.0472X0.1063*%
%ADD46O,0.0236X0.0472*%
%ADD47R,0.0591X0.0472*%
%ADD48R,0.0394X0.0374*%
%ADD49R,0.0374X0.0394*%
%ADD50R,0.1417X0.0551*%
%ADD51R,0.0866X0.0984*%
%ADD52R,0.0787X0.0197*%
%ADD53O,0.1062X0.0236*%
%ADD54O,0.0591X0.0256*%
%ADD55R,0.0197X0.0236*%
%ADD56R,0.0236X0.0197*%
%ADD57R,0.0236X0.0394*%
%ADD58R,0.0394X0.0236*%
%ADD59R,0.0236X0.0433*%
%ADD60R,0.0433X0.0236*%
%ADD61O,0.0571X0.0236*%
%ADD62O,0.0709X0.0591*%
%ADD63C,0.0708*%
%ADD64R,0.0708X0.0708*%
%ADD65R,0.0980X0.1370*%
%ADD66O,0.0591X0.0118*%
%ADD67R,0.0866X0.0630*%
%ADD68R,0.0177X0.0748*%
%ADD69O,0.0512X0.0236*%
%ADD70O,0.0866X0.0236*%
%ADD71R,0.1496X0.1496*%
%ADD72O,0.0118X0.0394*%
%ADD73O,0.0394X0.0118*%
%ADD74R,0.0472X0.0571*%
%ADD75R,0.1024X0.0945*%
%ADD76O,0.0118X0.0354*%
%ADD77O,0.0354X0.0118*%
%ADD78C,0.0394*%
%ADD79R,0.1969X0.1969*%
%ADD80R,0.0591X0.0118*%
%ADD81R,0.0118X0.0591*%
%ADD82R,0.0236X0.0453*%
%ADD83R,0.0453X0.0236*%
%ADD84R,0.0768X0.0866*%
%ADD85O,0.0630X0.0118*%
%ADD86R,0.0650X0.1949*%
%ADD87C,0.0197*%
%ADD88C,0.0394*%
%ADD89C,0.0118*%
%ADD90THERMAL90*%
%ADD91C,0.0787*%
%ADD92C,0.0630*%
%ADD93C,0.0550*%
%ADD94THERMAL94*%
%ADD95C,0.0709*%
%ADD96THERMAL96*%
%ADD97C,0.0709*%
%ADD98THERMAL98*%
%ADD99C,0.0591*%
%ADD100C,0.0866*%
%ADD101C,0.1378*%
%ADD102R,0.0709X0.0709*%
%ADD103C,0.1575*%
%ADD104O,0.1575X0.0787*%
%ADD105O,0.0787X0.1575*%
%ADD106O,0.0787X0.1772*%
%ADD107THERMAL107*%
%ADD108C,0.0709*%
%ADD109THERMAL109*%
%ADD110C,0.0709*%
%ADD111C,0.0050*%
%ADD112C,0.0050*%
%ADD113C,0.0315*%
%ADD114C,0.0050*%
%ADD115C,0.0050*%
%ADD116C,0.0315*%
%ADD117C,0.0217*%
%ADD118THERMAL118*%
%ADD119C,0.1181*%
%ADD120THERMAL120*%
%ADD121C,0.1181*%
%ADD122C,0.0750*%
%ADD123THERMAL123*%
%ADD124C,0.0217*%
%ADD125C,0.0217*%
%ADD126C,0.0050*%
%ADD127C,0.0217*%
%ADD128C,0.0050*%
%ADD129C,0.0787*%
%ADD130C,0.0630*%
%ADD131C,0.0550*%
%ADD132C,0.0709*%
%ADD133R,0.0709X0.0709*%
%ADD134C,0.0591*%
%ADD135THERMAL135*%
%ADD136R,0.0709X0.0709*%
%ADD137R,0.0709X0.0709*%
%ADD138C,0.0217*%
%ADD139THERMAL139*%
%ADD140C,0.1575*%
%ADD141C,0.0787*%
%ADD142C,0.0630*%
%ADD143C,0.0550*%
%ADD144C,0.0709*%
%ADD145R,0.0709X0.0709*%
%ADD146C,0.0591*%
%ADD147C,0.0866*%
%ADD148C,0.1378*%
%ADD149C,0.1575*%
%ADD150O,0.1575X0.0787*%
%ADD151O,0.0787X0.1575*%
%ADD152O,0.0787X0.1772*%
%ADD153C,0.0315*%
%ADD154C,0.0157*%
%ADD155C,0.0157*%
%ADD156C,0.0039*%
%ADD157R,0.0662X0.0583*%
%ADD158C,0.0004*%
%ADD159C,0.0157*%
%ADD160C,0.0000*%
%ADD161C,0.0078*%
%ADD162C,0.0100*%
%ADD163C,0.0020*%
%ADD164C,0.0071*%
%ADD165C,0.0067*%
%ADD166C,0.0070*%
%ADD167C,0.0059*%
*
G04 Plot Data ***
*
G54D29*
G01X0037491Y-0033021D02*
X0037403D01*
X0037447D02*
Y-0032758D01*
X0037403Y-0032802D01*
X0037158Y-0032889D02*
X0037180Y-0032846D01*
Y-0032802D01*
X0037158Y-0032758D01*
X0037027D01*
X0037005Y-0032802D01*
Y-0032846D01*
X0037027Y-0032889D01*
X0037158D01*
X0037180Y-0032933D01*
Y-0032977D01*
X0037158Y-0033021D01*
X0037027D01*
X0037005Y-0032977D01*
Y-0032933D01*
X0037027Y-0032889D01*
X0036826Y-0033021D02*
X0036739D01*
X0036782D02*
Y-0032758D01*
X0036739Y-0032802D01*
X0036516Y-0032758D02*
Y-0032846D01*
X0036428Y-0033021D01*
X0036341Y-0032846D01*
Y-0032758D01*
X0035986Y-0032889D02*
X0036117D01*
X0036161Y-0032846D01*
Y-0032802D01*
X0036117Y-0032758D01*
X0035986D01*
Y-0033021D01*
X0037425Y-0032509D02*
X0037381Y-0032465D01*
X0037359Y-0032421D01*
Y-0032334D01*
X0037381Y-0032290D01*
X0037425Y-0032246D01*
X0037469D01*
X0037513Y-0032290D01*
X0037535Y-0032334D01*
Y-0032421D01*
X0037513Y-0032465D01*
X0037469Y-0032509D01*
X0037425D01*
X0037158Y-0032378D02*
X0037180Y-0032334D01*
Y-0032290D01*
X0037158Y-0032246D01*
X0037027D01*
X0037005Y-0032290D01*
Y-0032334D01*
X0037027Y-0032378D01*
X0037158D01*
X0037180Y-0032421D01*
Y-0032465D01*
X0037158Y-0032509D01*
X0037027D01*
X0037005Y-0032465D01*
Y-0032421D01*
X0037027Y-0032378D01*
X0036826Y-0032509D02*
X0036739D01*
X0036782D02*
Y-0032246D01*
X0036739Y-0032290D01*
X0036516Y-0032246D02*
Y-0032334D01*
X0036428Y-0032509D01*
X0036341Y-0032334D01*
Y-0032246D01*
X0035986Y-0032378D02*
X0036117D01*
X0036161Y-0032334D01*
Y-0032290D01*
X0036117Y-0032246D01*
X0035986D01*
Y-0032509D01*
X0037513Y-0031866D02*
X0037381D01*
X0037359Y-0031822D01*
Y-0031778D01*
X0037381Y-0031735D01*
X0037513D01*
X0037535Y-0031778D01*
Y-0031822D01*
X0037447Y-0031997D01*
X0037049D02*
X0037180Y-0031735D01*
X0037005D01*
X0036826Y-0031997D02*
X0036739D01*
X0036782D02*
Y-0031735D01*
X0036739Y-0031778D01*
X0036516Y-0031735D02*
Y-0031822D01*
X0036428Y-0031997D01*
X0036341Y-0031822D01*
Y-0031735D01*
X0035986Y-0031866D02*
X0036117D01*
X0036161Y-0031822D01*
Y-0031778D01*
X0036117Y-0031735D01*
X0035986D01*
Y-0031997D01*
X0037001Y-0033913D02*
X0037023Y-0033869D01*
Y-0033826D01*
X0037001Y-0033782D01*
X0036870D01*
X0036848Y-0033826D01*
Y-0033869D01*
X0036870Y-0033913D01*
X0037001D01*
X0037023Y-0033957D01*
Y-0034001D01*
X0037001Y-0034044D01*
X0036870D01*
X0036848Y-0034001D01*
Y-0033957D01*
X0036870Y-0033913D01*
X0036537Y-0034044D02*
X0036669Y-0033782D01*
X0036493D01*
X0036314Y-0034044D02*
X0036227D01*
X0036270D02*
Y-0033782D01*
X0036227Y-0033826D01*
X0036004Y-0033782D02*
Y-0033869D01*
X0035916Y-0034044D01*
X0035829Y-0033869D01*
Y-0033782D01*
X0035474Y-0033913D02*
X0035606D01*
X0035650Y-0033869D01*
Y-0033826D01*
X0035606Y-0033782D01*
X0035474D01*
Y-0034044D01*
X0036891Y-0033533D02*
X0037023Y-0033270D01*
X0036848D01*
X0036537Y-0033533D02*
X0036669Y-0033270D01*
X0036493D01*
X0036314Y-0033533D02*
X0036227D01*
X0036270D02*
Y-0033270D01*
X0036227Y-0033314D01*
X0036004Y-0033270D02*
Y-0033357D01*
X0035916Y-0033533D01*
X0035829Y-0033357D01*
Y-0033270D01*
X0035474Y-0033401D02*
X0035606D01*
X0035650Y-0033357D01*
Y-0033314D01*
X0035606Y-0033270D01*
X0035474D01*
Y-0033533D01*
X0036870Y-0032889D02*
X0037001D01*
X0037023Y-0032933D01*
Y-0032977D01*
X0037001Y-0033021D01*
X0036870D01*
X0036848Y-0032977D01*
Y-0032933D01*
X0036935Y-0032758D01*
X0036537Y-0033021D02*
X0036669Y-0032758D01*
X0036493D01*
X0036314Y-0033021D02*
X0036227D01*
X0036270D02*
Y-0032758D01*
X0036227Y-0032802D01*
X0036004Y-0032758D02*
Y-0032846D01*
X0035916Y-0033021D01*
X0035829Y-0032846D01*
Y-0032758D01*
X0035474Y-0032889D02*
X0035606D01*
X0035650Y-0032846D01*
Y-0032802D01*
X0035606Y-0032758D01*
X0035474D01*
Y-0033021D01*
X0036848Y-0032465D02*
X0036870Y-0032509D01*
X0037001D01*
X0037023Y-0032465D01*
Y-0032378D01*
X0036979Y-0032334D01*
X0036848D01*
Y-0032246D01*
X0037023D01*
X0036537Y-0032509D02*
X0036669Y-0032246D01*
X0036493D01*
X0036314Y-0032509D02*
X0036227D01*
X0036270D02*
Y-0032246D01*
X0036227Y-0032290D01*
X0036004Y-0032246D02*
Y-0032334D01*
X0035916Y-0032509D01*
X0035829Y-0032334D01*
Y-0032246D01*
X0035474Y-0032378D02*
X0035606D01*
X0035650Y-0032334D01*
Y-0032290D01*
X0035606Y-0032246D01*
X0035474D01*
Y-0032509D01*
X0037023Y-0031909D02*
X0036848D01*
X0036935Y-0031735D01*
X0036979D01*
Y-0031997D01*
X0036537D02*
X0036669Y-0031735D01*
X0036493D01*
X0036314Y-0031997D02*
X0036227D01*
X0036270D02*
Y-0031735D01*
X0036227Y-0031778D01*
X0036004Y-0031735D02*
Y-0031822D01*
X0035916Y-0031997D01*
X0035829Y-0031822D01*
Y-0031735D01*
X0035474Y-0031866D02*
X0035606D01*
X0035650Y-0031822D01*
Y-0031778D01*
X0035606Y-0031735D01*
X0035474D01*
Y-0031997D01*
X0038383Y-0034001D02*
X0038427Y-0034044D01*
X0038514D01*
X0038558Y-0034001D01*
Y-0033957D01*
X0038470Y-0033869D01*
X0038558Y-0033782D01*
X0038383D01*
X0038182Y-0033913D02*
X0038051D01*
X0038029Y-0033869D01*
Y-0033826D01*
X0038051Y-0033782D01*
X0038182D01*
X0038204Y-0033826D01*
Y-0033869D01*
X0038116Y-0034044D01*
X0037850D02*
X0037762D01*
X0037806D02*
Y-0033782D01*
X0037762Y-0033826D01*
X0037539Y-0033782D02*
Y-0033869D01*
X0037452Y-0034044D01*
X0037364Y-0033869D01*
Y-0033782D01*
X0037010Y-0033913D02*
X0037141D01*
X0037185Y-0033869D01*
Y-0033826D01*
X0037141Y-0033782D01*
X0037010D01*
Y-0034044D01*
X0038558Y-0033533D02*
X0038383D01*
X0038558Y-0033357D01*
Y-0033314D01*
X0038536Y-0033270D01*
X0038405D01*
X0038383Y-0033314D01*
X0038182Y-0033401D02*
X0038051D01*
X0038029Y-0033357D01*
Y-0033314D01*
X0038051Y-0033270D01*
X0038182D01*
X0038204Y-0033314D01*
Y-0033357D01*
X0038116Y-0033533D01*
X0037850D02*
X0037762D01*
X0037806D02*
Y-0033270D01*
X0037762Y-0033314D01*
X0037539Y-0033270D02*
Y-0033357D01*
X0037452Y-0033533D01*
X0037364Y-0033357D01*
Y-0033270D01*
X0037010Y-0033401D02*
X0037141D01*
X0037185Y-0033357D01*
Y-0033314D01*
X0037141Y-0033270D01*
X0037010D01*
Y-0033533D01*
X0038514Y-0033021D02*
X0038427D01*
X0038470D02*
Y-0032758D01*
X0038427Y-0032802D01*
X0038182Y-0032889D02*
X0038051D01*
X0038029Y-0032846D01*
Y-0032802D01*
X0038051Y-0032758D01*
X0038182D01*
X0038204Y-0032802D01*
Y-0032846D01*
X0038116Y-0033021D01*
X0037850D02*
X0037762D01*
X0037806D02*
Y-0032758D01*
X0037762Y-0032802D01*
X0037539Y-0032758D02*
Y-0032846D01*
X0037452Y-0033021D01*
X0037364Y-0032846D01*
Y-0032758D01*
X0037010Y-0032889D02*
X0037141D01*
X0037185Y-0032846D01*
Y-0032802D01*
X0037141Y-0032758D01*
X0037010D01*
Y-0033021D01*
X0038449Y-0032509D02*
X0038405Y-0032465D01*
X0038383Y-0032421D01*
Y-0032334D01*
X0038405Y-0032290D01*
X0038449Y-0032246D01*
X0038493D01*
X0038536Y-0032290D01*
X0038558Y-0032334D01*
Y-0032421D01*
X0038536Y-0032465D01*
X0038493Y-0032509D01*
X0038449D01*
X0038182Y-0032378D02*
X0038051D01*
X0038029Y-0032334D01*
Y-0032290D01*
X0038051Y-0032246D01*
X0038182D01*
X0038204Y-0032290D01*
Y-0032334D01*
X0038116Y-0032509D01*
X0037850D02*
X0037762D01*
X0037806D02*
Y-0032246D01*
X0037762Y-0032290D01*
X0037539Y-0032246D02*
Y-0032334D01*
X0037452Y-0032509D01*
X0037364Y-0032334D01*
Y-0032246D01*
X0037010Y-0032378D02*
X0037141D01*
X0037185Y-0032334D01*
Y-0032290D01*
X0037141Y-0032246D01*
X0037010D01*
Y-0032509D01*
X0038536Y-0031866D02*
X0038405D01*
X0038383Y-0031822D01*
Y-0031778D01*
X0038405Y-0031735D01*
X0038536D01*
X0038558Y-0031778D01*
Y-0031822D01*
X0038470Y-0031997D01*
X0038182Y-0031866D02*
X0038204Y-0031822D01*
Y-0031778D01*
X0038182Y-0031735D01*
X0038051D01*
X0038029Y-0031778D01*
Y-0031822D01*
X0038051Y-0031866D01*
X0038182D01*
X0038204Y-0031909D01*
Y-0031954D01*
X0038182Y-0031997D01*
X0038051D01*
X0038029Y-0031954D01*
Y-0031909D01*
X0038051Y-0031866D01*
X0037850Y-0031997D02*
X0037762D01*
X0037806D02*
Y-0031735D01*
X0037762Y-0031778D01*
X0037539Y-0031735D02*
Y-0031822D01*
X0037452Y-0031997D01*
X0037364Y-0031822D01*
Y-0031735D01*
X0037010Y-0031866D02*
X0037141D01*
X0037185Y-0031822D01*
Y-0031778D01*
X0037141Y-0031735D01*
X0037010D01*
Y-0031997D01*
X0038024Y-0033401D02*
X0038046Y-0033357D01*
Y-0033314D01*
X0038024Y-0033270D01*
X0037893D01*
X0037871Y-0033314D01*
Y-0033357D01*
X0037893Y-0033401D01*
X0038024D01*
X0038046Y-0033445D01*
Y-0033489D01*
X0038024Y-0033533D01*
X0037893D01*
X0037871Y-0033489D01*
Y-0033445D01*
X0037893Y-0033401D01*
X0037670D02*
X0037692Y-0033357D01*
Y-0033314D01*
X0037670Y-0033270D01*
X0037539D01*
X0037517Y-0033314D01*
Y-0033357D01*
X0037539Y-0033401D01*
X0037670D01*
X0037692Y-0033445D01*
Y-0033489D01*
X0037670Y-0033533D01*
X0037539D01*
X0037517Y-0033489D01*
Y-0033445D01*
X0037539Y-0033401D01*
X0037338Y-0033533D02*
X0037250D01*
X0037294D02*
Y-0033270D01*
X0037250Y-0033314D01*
X0037028Y-0033270D02*
Y-0033357D01*
X0036940Y-0033533D01*
X0036852Y-0033357D01*
Y-0033270D01*
X0036498Y-0033401D02*
X0036629D01*
X0036673Y-0033357D01*
Y-0033314D01*
X0036629Y-0033270D01*
X0036498D01*
Y-0033533D01*
X0037915Y-0033021D02*
X0038046Y-0032758D01*
X0037871D01*
X0037670Y-0032889D02*
X0037692Y-0032846D01*
Y-0032802D01*
X0037670Y-0032758D01*
X0037539D01*
X0037517Y-0032802D01*
Y-0032846D01*
X0037539Y-0032889D01*
X0037670D01*
X0037692Y-0032933D01*
Y-0032977D01*
X0037670Y-0033021D01*
X0037539D01*
X0037517Y-0032977D01*
Y-0032933D01*
X0037539Y-0032889D01*
X0037338Y-0033021D02*
X0037250D01*
X0037294D02*
Y-0032758D01*
X0037250Y-0032802D01*
X0037028Y-0032758D02*
Y-0032846D01*
X0036940Y-0033021D01*
X0036852Y-0032846D01*
Y-0032758D01*
X0036498Y-0032889D02*
X0036629D01*
X0036673Y-0032846D01*
Y-0032802D01*
X0036629Y-0032758D01*
X0036498D01*
Y-0033021D01*
X0037893Y-0032378D02*
X0038024D01*
X0038046Y-0032421D01*
Y-0032465D01*
X0038024Y-0032509D01*
X0037893D01*
X0037871Y-0032465D01*
Y-0032421D01*
X0037959Y-0032246D01*
X0037670Y-0032378D02*
X0037692Y-0032334D01*
Y-0032290D01*
X0037670Y-0032246D01*
X0037539D01*
X0037517Y-0032290D01*
Y-0032334D01*
X0037539Y-0032378D01*
X0037670D01*
X0037692Y-0032421D01*
Y-0032465D01*
X0037670Y-0032509D01*
X0037539D01*
X0037517Y-0032465D01*
Y-0032421D01*
X0037539Y-0032378D01*
X0037338Y-0032509D02*
X0037250D01*
X0037294D02*
Y-0032246D01*
X0037250Y-0032290D01*
X0037028Y-0032246D02*
Y-0032334D01*
X0036940Y-0032509D01*
X0036852Y-0032334D01*
Y-0032246D01*
X0036498Y-0032378D02*
X0036629D01*
X0036673Y-0032334D01*
Y-0032290D01*
X0036629Y-0032246D01*
X0036498D01*
Y-0032509D01*
X0037871Y-0031954D02*
X0037893Y-0031997D01*
X0038024D01*
X0038046Y-0031954D01*
Y-0031866D01*
X0038002Y-0031822D01*
X0037871D01*
Y-0031735D01*
X0038046D01*
X0037670Y-0031866D02*
X0037692Y-0031822D01*
Y-0031778D01*
X0037670Y-0031735D01*
X0037539D01*
X0037517Y-0031778D01*
Y-0031822D01*
X0037539Y-0031866D01*
X0037670D01*
X0037692Y-0031909D01*
Y-0031954D01*
X0037670Y-0031997D01*
X0037539D01*
X0037517Y-0031954D01*
Y-0031909D01*
X0037539Y-0031866D01*
X0037338Y-0031997D02*
X0037250D01*
X0037294D02*
Y-0031735D01*
X0037250Y-0031778D01*
X0037028Y-0031735D02*
Y-0031822D01*
X0036940Y-0031997D01*
X0036852Y-0031822D01*
Y-0031735D01*
X0036498Y-0031866D02*
X0036629D01*
X0036673Y-0031822D01*
Y-0031778D01*
X0036629Y-0031735D01*
X0036498D01*
Y-0031997D01*
X0038046Y-0033957D02*
X0037871D01*
X0037959Y-0033782D01*
X0038002D01*
Y-0034044D01*
X0037670Y-0033913D02*
X0037692Y-0033869D01*
Y-0033826D01*
X0037670Y-0033782D01*
X0037539D01*
X0037517Y-0033826D01*
Y-0033869D01*
X0037539Y-0033913D01*
X0037670D01*
X0037692Y-0033957D01*
Y-0034001D01*
X0037670Y-0034044D01*
X0037539D01*
X0037517Y-0034001D01*
Y-0033957D01*
X0037539Y-0033913D01*
X0037338Y-0034044D02*
X0037250D01*
X0037294D02*
Y-0033782D01*
X0037250Y-0033826D01*
X0037028Y-0033782D02*
Y-0033869D01*
X0036940Y-0034044D01*
X0036852Y-0033869D01*
Y-0033782D01*
X0036498Y-0033913D02*
X0036629D01*
X0036673Y-0033869D01*
Y-0033826D01*
X0036629Y-0033782D01*
X0036498D01*
Y-0034044D01*
X0037359Y-0034001D02*
X0037403Y-0034044D01*
X0037491D01*
X0037535Y-0034001D01*
Y-0033957D01*
X0037447Y-0033869D01*
X0037535Y-0033782D01*
X0037359D01*
X0037158Y-0033913D02*
X0037180Y-0033869D01*
Y-0033826D01*
X0037158Y-0033782D01*
X0037027D01*
X0037005Y-0033826D01*
Y-0033869D01*
X0037027Y-0033913D01*
X0037158D01*
X0037180Y-0033957D01*
Y-0034001D01*
X0037158Y-0034044D01*
X0037027D01*
X0037005Y-0034001D01*
Y-0033957D01*
X0037027Y-0033913D01*
X0036826Y-0034044D02*
X0036739D01*
X0036782D02*
Y-0033782D01*
X0036739Y-0033826D01*
X0036516Y-0033782D02*
Y-0033869D01*
X0036428Y-0034044D01*
X0036341Y-0033869D01*
Y-0033782D01*
X0035986Y-0033913D02*
X0036117D01*
X0036161Y-0033869D01*
Y-0033826D01*
X0036117Y-0033782D01*
X0035986D01*
Y-0034044D01*
X0037535Y-0033533D02*
X0037359D01*
X0037535Y-0033357D01*
Y-0033314D01*
X0037513Y-0033270D01*
X0037381D01*
X0037359Y-0033314D01*
X0037158Y-0033401D02*
X0037180Y-0033357D01*
Y-0033314D01*
X0037158Y-0033270D01*
X0037027D01*
X0037005Y-0033314D01*
Y-0033357D01*
X0037027Y-0033401D01*
X0037158D01*
X0037180Y-0033445D01*
Y-0033489D01*
X0037158Y-0033533D01*
X0037027D01*
X0037005Y-0033489D01*
Y-0033445D01*
X0037027Y-0033401D01*
X0036826Y-0033533D02*
X0036739D01*
X0036782D02*
Y-0033270D01*
X0036739Y-0033314D01*
X0036516Y-0033270D02*
Y-0033357D01*
X0036428Y-0033533D01*
X0036341Y-0033357D01*
Y-0033270D01*
X0035986Y-0033401D02*
X0036117D01*
X0036161Y-0033357D01*
Y-0033314D01*
X0036117Y-0033270D01*
X0035986D01*
Y-0033533D01*
X0038335Y-0034110D02*
X0038357Y-0034066D01*
Y-0034022D01*
X0038335Y-0033979D01*
X0038204D01*
X0038181Y-0034022D01*
Y-0034066D01*
X0038204Y-0034110D01*
X0038335D01*
X0038357Y-0034154D01*
Y-0034198D01*
X0038335Y-0034241D01*
X0038204D01*
X0038181Y-0034198D01*
Y-0034154D01*
X0038204Y-0034110D01*
X0038002Y-0034241D02*
X0037915D01*
X0037959D02*
Y-0033979D01*
X0037915Y-0034022D01*
X0037692Y-0034241D02*
X0037605D01*
X0037648D02*
Y-0033979D01*
X0037605Y-0034022D01*
X0037382Y-0033979D02*
Y-0034066D01*
X0037294Y-0034241D01*
X0037207Y-0034066D01*
Y-0033979D01*
X0036852Y-0034110D02*
X0036983D01*
X0037028Y-0034066D01*
Y-0034022D01*
X0036983Y-0033979D01*
X0036852D01*
Y-0034241D01*
X0038225Y-0033730D02*
X0038357Y-0033467D01*
X0038181D01*
X0038002Y-0033730D02*
X0037915D01*
X0037959D02*
Y-0033467D01*
X0037915Y-0033511D01*
X0037692Y-0033730D02*
X0037605D01*
X0037648D02*
Y-0033467D01*
X0037605Y-0033511D01*
X0037382Y-0033467D02*
Y-0033554D01*
X0037294Y-0033730D01*
X0037207Y-0033554D01*
Y-0033467D01*
X0036852Y-0033598D02*
X0036983D01*
X0037028Y-0033554D01*
Y-0033511D01*
X0036983Y-0033467D01*
X0036852D01*
Y-0033730D01*
X0037180Y-0033598D02*
X0037311D01*
X0037333Y-0033642D01*
Y-0033686D01*
X0037311Y-0033730D01*
X0037180D01*
X0037158Y-0033686D01*
Y-0033642D01*
X0037245Y-0033467D01*
X0036979Y-0033730D02*
X0036891D01*
X0036935D02*
Y-0033467D01*
X0036891Y-0033511D01*
X0036669Y-0033730D02*
X0036581D01*
X0036625D02*
Y-0033467D01*
X0036581Y-0033511D01*
X0036358Y-0033467D02*
Y-0033554D01*
X0036270Y-0033730D01*
X0036183Y-0033554D01*
Y-0033467D01*
X0035829Y-0033598D02*
X0035960D01*
X0036004Y-0033554D01*
Y-0033511D01*
X0035960Y-0033467D01*
X0035829D01*
Y-0033730D01*
X0036646Y-0032150D02*
X0036668Y-0032194D01*
X0036799D01*
X0036821Y-0032150D01*
Y-0032063D01*
X0036777Y-0032019D01*
X0036646D01*
Y-0031931D01*
X0036821D01*
X0036467Y-0032194D02*
X0036380D01*
X0036423D02*
Y-0031931D01*
X0036380Y-0031975D01*
X0036157Y-0032194D02*
X0036069D01*
X0036113D02*
Y-0031931D01*
X0036069Y-0031975D01*
X0035846Y-0031931D02*
Y-0032019D01*
X0035759Y-0032194D01*
X0035671Y-0032019D01*
Y-0031931D01*
X0035317Y-0032063D02*
X0035448D01*
X0035492Y-0032019D01*
Y-0031975D01*
X0035448Y-0031931D01*
X0035317D01*
Y-0032194D01*
X0036821Y-0033642D02*
X0036646D01*
X0036733Y-0033467D01*
X0036777D01*
Y-0033730D01*
X0036467D02*
X0036380D01*
X0036423D02*
Y-0033467D01*
X0036380Y-0033511D01*
X0036157Y-0033730D02*
X0036069D01*
X0036113D02*
Y-0033467D01*
X0036069Y-0033511D01*
X0035846Y-0033467D02*
Y-0033554D01*
X0035759Y-0033730D01*
X0035671Y-0033554D01*
Y-0033467D01*
X0035317Y-0033598D02*
X0035448D01*
X0035492Y-0033554D01*
Y-0033511D01*
X0035448Y-0033467D01*
X0035317D01*
Y-0033730D01*
X0037670Y-0034198D02*
X0037713Y-0034241D01*
X0037801D01*
X0037845Y-0034198D01*
Y-0034154D01*
X0037757Y-0034066D01*
X0037845Y-0033979D01*
X0037670D01*
X0037491Y-0034241D02*
X0037403D01*
X0037447D02*
Y-0033979D01*
X0037403Y-0034022D01*
X0037180Y-0034241D02*
X0037093D01*
X0037137D02*
Y-0033979D01*
X0037093Y-0034022D01*
X0036870Y-0033979D02*
Y-0034066D01*
X0036782Y-0034241D01*
X0036695Y-0034066D01*
Y-0033979D01*
X0036341Y-0034110D02*
X0036472D01*
X0036516Y-0034066D01*
Y-0034022D01*
X0036472Y-0033979D01*
X0036341D01*
Y-0034241D01*
X0037845Y-0033730D02*
X0037670D01*
X0037845Y-0033554D01*
Y-0033511D01*
X0037823Y-0033467D01*
X0037692D01*
X0037670Y-0033511D01*
X0037491Y-0033730D02*
X0037403D01*
X0037447D02*
Y-0033467D01*
X0037403Y-0033511D01*
X0037180Y-0033730D02*
X0037093D01*
X0037137D02*
Y-0033467D01*
X0037093Y-0033511D01*
X0036870Y-0033467D02*
Y-0033554D01*
X0036782Y-0033730D01*
X0036695Y-0033554D01*
Y-0033467D01*
X0036341Y-0033598D02*
X0036472D01*
X0036516Y-0033554D01*
Y-0033511D01*
X0036472Y-0033467D01*
X0036341D01*
Y-0033730D01*
X0036690Y-0033174D02*
X0036712Y-0033218D01*
X0036843D01*
X0036865Y-0033174D01*
Y-0033086D01*
X0036821Y-0033043D01*
X0036690D01*
Y-0032955D01*
X0036865D01*
X0036358Y-0033086D02*
X0036489D01*
X0036511Y-0033130D01*
Y-0033174D01*
X0036489Y-0033218D01*
X0036358D01*
X0036336Y-0033174D01*
Y-0033130D01*
X0036423Y-0032955D01*
X0036157Y-0033218D02*
X0036069D01*
X0036113D02*
Y-0032955D01*
X0036069Y-0032999D01*
X0035846Y-0032955D02*
Y-0033043D01*
X0035759Y-0033218D01*
X0035671Y-0033043D01*
Y-0032955D01*
X0035317Y-0033086D02*
X0035448D01*
X0035492Y-0033043D01*
Y-0032999D01*
X0035448Y-0032955D01*
X0035317D01*
Y-0033218D01*
X0038401Y-0033130D02*
X0038226D01*
X0038313Y-0032955D01*
X0038357D01*
Y-0033218D01*
X0037893Y-0033086D02*
X0038024D01*
X0038046Y-0033130D01*
Y-0033174D01*
X0038024Y-0033218D01*
X0037893D01*
X0037871Y-0033174D01*
Y-0033130D01*
X0037959Y-0032955D01*
X0037692Y-0033218D02*
X0037605D01*
X0037648D02*
Y-0032955D01*
X0037605Y-0032999D01*
X0037382Y-0032955D02*
Y-0033043D01*
X0037294Y-0033218D01*
X0037207Y-0033043D01*
Y-0032955D01*
X0036852Y-0033086D02*
X0036983D01*
X0037028Y-0033043D01*
Y-0032999D01*
X0036983Y-0032955D01*
X0036852D01*
Y-0033218D01*
X0037714Y-0032662D02*
X0037757Y-0032706D01*
X0037845D01*
X0037889Y-0032662D01*
Y-0032618D01*
X0037801Y-0032531D01*
X0037889Y-0032443D01*
X0037714D01*
X0037381Y-0032574D02*
X0037513D01*
X0037535Y-0032618D01*
Y-0032662D01*
X0037513Y-0032706D01*
X0037381D01*
X0037359Y-0032662D01*
Y-0032618D01*
X0037447Y-0032443D01*
X0037180Y-0032706D02*
X0037093D01*
X0037137D02*
Y-0032443D01*
X0037093Y-0032487D01*
X0036870Y-0032443D02*
Y-0032531D01*
X0036782Y-0032706D01*
X0036695Y-0032531D01*
Y-0032443D01*
X0036341Y-0032574D02*
X0036472D01*
X0036516Y-0032531D01*
Y-0032487D01*
X0036472Y-0032443D01*
X0036341D01*
Y-0032706D01*
X0037377D02*
X0037202D01*
X0037377Y-0032531D01*
Y-0032487D01*
X0037355Y-0032443D01*
X0037224D01*
X0037202Y-0032487D01*
X0036870Y-0032574D02*
X0037001D01*
X0037023Y-0032618D01*
Y-0032662D01*
X0037001Y-0032706D01*
X0036870D01*
X0036848Y-0032662D01*
Y-0032618D01*
X0036935Y-0032443D01*
X0036669Y-0032706D02*
X0036581D01*
X0036625D02*
Y-0032443D01*
X0036581Y-0032487D01*
X0036358Y-0032443D02*
Y-0032531D01*
X0036270Y-0032706D01*
X0036183Y-0032531D01*
Y-0032443D01*
X0035829Y-0032574D02*
X0035960D01*
X0036004Y-0032531D01*
Y-0032487D01*
X0035960Y-0032443D01*
X0035829D01*
Y-0032706D01*
X0037355Y-0032063D02*
X0037224D01*
X0037202Y-0032019D01*
Y-0031975D01*
X0037224Y-0031931D01*
X0037355D01*
X0037377Y-0031975D01*
Y-0032019D01*
X0037289Y-0032194D01*
X0036870Y-0032063D02*
X0037001D01*
X0037023Y-0032106D01*
Y-0032150D01*
X0037001Y-0032194D01*
X0036870D01*
X0036848Y-0032150D01*
Y-0032106D01*
X0036935Y-0031931D01*
X0036669Y-0032194D02*
X0036581D01*
X0036625D02*
Y-0031931D01*
X0036581Y-0031975D01*
X0036358Y-0031931D02*
Y-0032019D01*
X0036270Y-0032194D01*
X0036183Y-0032019D01*
Y-0031931D01*
X0035829Y-0032063D02*
X0035960D01*
X0036004Y-0032019D01*
Y-0031975D01*
X0035960Y-0031931D01*
X0035829D01*
Y-0032194D01*
X0038379Y-0032574D02*
X0038401Y-0032531D01*
Y-0032487D01*
X0038379Y-0032443D01*
X0038248D01*
X0038226Y-0032487D01*
Y-0032531D01*
X0038248Y-0032574D01*
X0038379D01*
X0038401Y-0032618D01*
Y-0032662D01*
X0038379Y-0032706D01*
X0038248D01*
X0038226Y-0032662D01*
Y-0032618D01*
X0038248Y-0032574D01*
X0037893D02*
X0038024D01*
X0038046Y-0032618D01*
Y-0032662D01*
X0038024Y-0032706D01*
X0037893D01*
X0037871Y-0032662D01*
Y-0032618D01*
X0037959Y-0032443D01*
X0037692Y-0032706D02*
X0037605D01*
X0037648D02*
Y-0032443D01*
X0037605Y-0032487D01*
X0037382Y-0032443D02*
Y-0032531D01*
X0037294Y-0032706D01*
X0037207Y-0032531D01*
Y-0032443D01*
X0036852Y-0032574D02*
X0036983D01*
X0037028Y-0032531D01*
Y-0032487D01*
X0036983Y-0032443D01*
X0036852D01*
Y-0032706D01*
X0037757Y-0033218D02*
X0037889Y-0032955D01*
X0037714D01*
X0037381Y-0033086D02*
X0037513D01*
X0037535Y-0033130D01*
Y-0033174D01*
X0037513Y-0033218D01*
X0037381D01*
X0037359Y-0033174D01*
Y-0033130D01*
X0037447Y-0032955D01*
X0037180Y-0033218D02*
X0037093D01*
X0037137D02*
Y-0032955D01*
X0037093Y-0032999D01*
X0036870Y-0032955D02*
Y-0033043D01*
X0036782Y-0033218D01*
X0036695Y-0033043D01*
Y-0032955D01*
X0036341Y-0033086D02*
X0036472D01*
X0036516Y-0033043D01*
Y-0032999D01*
X0036472Y-0032955D01*
X0036341D01*
Y-0033218D01*
X0036712Y-0032574D02*
X0036843D01*
X0036865Y-0032618D01*
Y-0032662D01*
X0036843Y-0032706D01*
X0036712D01*
X0036690Y-0032662D01*
Y-0032618D01*
X0036778Y-0032443D01*
X0036358Y-0032574D02*
X0036489D01*
X0036511Y-0032618D01*
Y-0032662D01*
X0036489Y-0032706D01*
X0036358D01*
X0036336Y-0032662D01*
Y-0032618D01*
X0036423Y-0032443D01*
X0036157Y-0032706D02*
X0036069D01*
X0036113D02*
Y-0032443D01*
X0036069Y-0032487D01*
X0035846Y-0032443D02*
Y-0032531D01*
X0035759Y-0032706D01*
X0035671Y-0032531D01*
Y-0032443D01*
X0035317Y-0032574D02*
X0035448D01*
X0035492Y-0032531D01*
Y-0032487D01*
X0035448Y-0032443D01*
X0035317D01*
Y-0032706D01*
X0037953Y0036620D02*
X0037909Y0036708D01*
X0037646D01*
X0037603Y0036620D01*
Y0036533D01*
X0037646Y0036446D01*
X0037909D01*
X0037953Y0036358D01*
Y0036270D01*
X0037909Y0036183D01*
X0037646D01*
X0037603Y0036270D01*
X0037270Y0036446D02*
X0037402Y0036183D01*
X0037052Y0036446D02*
X0037314D01*
X0037402Y0036533D01*
Y0036620D01*
X0037314Y0036708D01*
X0037052D01*
Y0036183D01*
X0036544D02*
X0036500Y0036270D01*
Y0036620D01*
X0036544Y0036708D01*
X0036806D01*
X0036850Y0036620D01*
Y0036270D01*
X0036806Y0036183D01*
X0036544D01*
X0036168Y0036446D02*
X0036299Y0036183D01*
X0035949Y0036446D02*
X0036211D01*
X0036299Y0036533D01*
Y0036620D01*
X0036211Y0036708D01*
X0035949D01*
Y0036183D01*
X0035617Y0036446D02*
X0035748Y0036183D01*
X0035398Y0036446D02*
X0035660D01*
X0035748Y0036533D01*
Y0036620D01*
X0035660Y0036708D01*
X0035398D01*
Y0036183D01*
X0035109Y0036446D02*
X0034847D01*
X0035197Y0036183D02*
X0034847D01*
Y0036708D01*
X0035197D01*
X0033591Y0036183D02*
Y0036708D01*
X0033548Y0036183D02*
X0033810D01*
X0033898Y0036358D01*
Y0036533D01*
X0033810Y0036708D01*
X0033548D01*
X0033040Y0036183D02*
X0032996Y0036270D01*
Y0036620D01*
X0033040Y0036708D01*
X0033302D01*
X0033346Y0036620D01*
Y0036270D01*
X0033302Y0036183D01*
X0033040D01*
X0032489D02*
X0032445Y0036270D01*
Y0036620D01*
X0032489Y0036708D01*
X0032751D01*
X0032795Y0036620D01*
Y0036270D01*
X0032751Y0036183D01*
X0032489D01*
X0032069Y0036446D02*
X0032244D01*
Y0036270D01*
X0032200Y0036183D01*
X0031938D01*
X0031894Y0036270D01*
Y0036620D01*
X0031938Y0036708D01*
X0032200D01*
X0032244Y0036620D01*
X0030945Y0036708D02*
Y0036183D01*
X0030857Y0036270D01*
X0030682Y0036620D01*
X0030595Y0036708D01*
Y0036183D01*
X0030394Y0036708D02*
Y0036270D01*
X0030350Y0036183D01*
X0030219Y0036446D01*
Y0036533D02*
Y0036446D01*
X0030087Y0036183D01*
X0030044Y0036270D01*
Y0036708D01*
X0029536Y0036183D02*
X0029493Y0036270D01*
Y0036620D01*
X0029536Y0036708D01*
X0029798D01*
X0029843Y0036620D01*
Y0036270D01*
X0029798Y0036183D01*
X0029536D01*
X0029291Y0036708D02*
Y0036183D01*
X0029204Y0036270D01*
X0029029Y0036620D01*
X0028941Y0036708D01*
Y0036183D01*
X0028740D02*
X0028478Y0036446D01*
X0028740Y0036708D01*
X0028390D02*
Y0036183D01*
X0027397Y0036446D02*
X0027441Y0036533D01*
Y0036620D01*
X0027397Y0036708D01*
X0027135D01*
X0027091Y0036620D01*
Y0036533D01*
X0027135Y0036446D01*
X0027397D01*
X0027441Y0036358D01*
Y0036270D01*
X0027397Y0036183D01*
X0027135D01*
X0027091Y0036270D01*
Y0036358D01*
X0027135Y0036446D01*
X0026890Y0036358D02*
X0026540D01*
X0026715Y0036708D01*
X0026802D01*
Y0036183D01*
X0031808Y-0032131D02*
X0031830Y-0032174D01*
X0031961D01*
X0031983Y-0032131D01*
Y-0032043D01*
X0031939Y-0031999D01*
X0031808D01*
Y-0031912D01*
X0031983D01*
X0031629Y-0032087D02*
X0031454D01*
X0031541Y-0031912D01*
X0031585D01*
Y-0032174D01*
X0031275D02*
X0031187D01*
X0031231D02*
Y-0031912D01*
X0031187Y-0031956D01*
X0030965Y-0031912D02*
Y-0031999D01*
X0030877Y-0032174D01*
X0030789Y-0031999D01*
Y-0031912D01*
X0030435Y-0032043D02*
X0030566D01*
X0030610Y-0031999D01*
Y-0031956D01*
X0030566Y-0031912D01*
X0030435D01*
Y-0032174D01*
X0032419Y-0031481D02*
X0032462Y-0031525D01*
X0032550D01*
X0032594Y-0031481D01*
Y-0031437D01*
X0032506Y-0031350D01*
X0032594Y-0031262D01*
X0032419D01*
X0032239Y-0031437D02*
X0032064D01*
X0032152Y-0031262D01*
X0032195D01*
Y-0031525D01*
X0031885D02*
X0031798D01*
X0031841D02*
Y-0031262D01*
X0031798Y-0031306D01*
X0031575Y-0031262D02*
Y-0031350D01*
X0031487Y-0031525D01*
X0031400Y-0031350D01*
Y-0031262D01*
X0031045Y-0031393D02*
X0031176D01*
X0031220Y-0031350D01*
Y-0031306D01*
X0031176Y-0031262D01*
X0031045D01*
Y-0031525D01*
X0037845Y-0032194D02*
X0037757D01*
X0037801D02*
Y-0031931D01*
X0037757Y-0031975D01*
X0037381Y-0032063D02*
X0037513D01*
X0037535Y-0032106D01*
Y-0032150D01*
X0037513Y-0032194D01*
X0037381D01*
X0037359Y-0032150D01*
Y-0032106D01*
X0037447Y-0031931D01*
X0037180Y-0032194D02*
X0037093D01*
X0037137D02*
Y-0031931D01*
X0037093Y-0031975D01*
X0036870Y-0031931D02*
Y-0032019D01*
X0036782Y-0032194D01*
X0036695Y-0032019D01*
Y-0031931D01*
X0036341Y-0032063D02*
X0036472D01*
X0036516Y-0032019D01*
Y-0031975D01*
X0036472Y-0031931D01*
X0036341D01*
Y-0032194D01*
X0037268Y-0033218D02*
X0037224Y-0033174D01*
X0037202Y-0033130D01*
Y-0033043D01*
X0037224Y-0032999D01*
X0037268Y-0032955D01*
X0037311D01*
X0037355Y-0032999D01*
X0037377Y-0033043D01*
Y-0033130D01*
X0037355Y-0033174D01*
X0037311Y-0033218D01*
X0037268D01*
X0036870Y-0033086D02*
X0037001D01*
X0037023Y-0033130D01*
Y-0033174D01*
X0037001Y-0033218D01*
X0036870D01*
X0036848Y-0033174D01*
Y-0033130D01*
X0036935Y-0032955D01*
X0036669Y-0033218D02*
X0036581D01*
X0036625D02*
Y-0032955D01*
X0036581Y-0032999D01*
X0036358Y-0032955D02*
Y-0033043D01*
X0036270Y-0033218D01*
X0036183Y-0033043D01*
Y-0032955D01*
X0035829Y-0033086D02*
X0035960D01*
X0036004Y-0033043D01*
Y-0032999D01*
X0035960Y-0032955D01*
X0035829D01*
Y-0033218D01*
X-0006687Y-0034812D02*
X-0006643Y-0034856D01*
X-0006556D01*
X-0006512Y-0034812D01*
Y-0034768D01*
X-0006600Y-0034680D01*
X-0006512Y-0034593D01*
X-0006687D01*
X-0007019Y-0034856D02*
Y-0034593D01*
X-0007041Y-0034856D02*
X-0006910D01*
X-0006866Y-0034768D01*
Y-0034680D01*
X-0006910Y-0034593D01*
X-0007041D01*
X-0007220Y-0034724D02*
X-0007396D01*
X-0007220Y-0034856D02*
Y-0034593D01*
X-0007396Y-0034856D02*
Y-0034593D01*
X-0019788Y0004311D02*
X-0019963D01*
X-0019876Y0004486D01*
X-0019832D01*
Y0004223D01*
X-0020143D02*
X-0020230D01*
X-0020186D02*
Y0004486D01*
X-0020230Y0004442D01*
X-0020453Y0004486D02*
Y0004267D01*
X-0020475Y0004223D01*
X-0020606D01*
X-0020628Y0004267D01*
Y0004486D01*
X0031983Y-0031437D02*
X0031808D01*
X0031896Y-0031262D01*
X0031939D01*
Y-0031525D01*
X0031629Y-0031437D02*
X0031454D01*
X0031541Y-0031262D01*
X0031585D01*
Y-0031525D01*
X0031275D02*
X0031187D01*
X0031231D02*
Y-0031262D01*
X0031187Y-0031306D01*
X0030965Y-0031262D02*
Y-0031350D01*
X0030877Y-0031525D01*
X0030789Y-0031350D01*
Y-0031262D01*
X0030435Y-0031393D02*
X0030566D01*
X0030610Y-0031350D01*
Y-0031306D01*
X0030566Y-0031262D01*
X0030435D01*
Y-0031525D01*
X0035089Y-0032740D02*
X0035133Y-0032696D01*
X0035177Y-0032674D01*
X0035265D01*
X0035308Y-0032696D01*
X0035352Y-0032740D01*
Y-0032784D01*
X0035308Y-0032828D01*
X0035265Y-0032850D01*
X0035177D01*
X0035133Y-0032828D01*
X0035089Y-0032784D01*
Y-0032740D01*
Y-0032495D02*
Y-0032408D01*
Y-0032452D02*
X0035352D01*
X0035308Y-0032408D01*
X0035352Y-0032185D02*
X0035265D01*
X0035089Y-0032097D01*
X0035265Y-0032010D01*
X0035352D01*
X0035221Y-0031656D02*
Y-0031787D01*
X0035265Y-0031831D01*
X0035308D01*
X0035352Y-0031787D01*
Y-0031656D01*
X0035089D01*
X-0005742Y0005345D02*
X-0005785Y0005389D01*
X-0005807Y0005433D01*
Y0005520D01*
X-0005785Y0005564D01*
X-0005742Y0005608D01*
X-0005698D01*
X-0005654Y0005564D01*
X-0005632Y0005520D01*
Y0005433D01*
X-0005654Y0005389D01*
X-0005698Y0005345D01*
X-0005742D01*
X-0006162Y0005389D02*
X-0006118Y0005345D01*
X-0006031D01*
X-0005987Y0005389D01*
Y0005433D01*
X-0006074Y0005520D01*
X-0005987Y0005608D01*
X-0006162D01*
X-0006494Y0005345D02*
Y0005608D01*
X-0006516Y0005345D02*
X-0006385D01*
X-0006341Y0005433D01*
Y0005520D01*
X-0006385Y0005608D01*
X-0006516D01*
X-0006739Y0005477D02*
X-0006870D01*
X-0006695Y0005345D02*
X-0006870D01*
Y0005608D01*
X-0006695D01*
X-0007050Y0005345D02*
X-0007203D01*
Y0005608D01*
X-0003922Y0005477D02*
X-0004053D01*
X-0004075Y0005520D01*
Y0005564D01*
X-0004053Y0005608D01*
X-0003922D01*
X-0003900Y0005564D01*
Y0005520D01*
X-0003988Y0005345D01*
X-0004254D02*
X-0004430D01*
X-0004254Y0005520D01*
Y0005564D01*
X-0004276Y0005608D01*
X-0004407D01*
X-0004430Y0005564D01*
X-0004762Y0005345D02*
Y0005608D01*
X-0004784Y0005345D02*
X-0004653D01*
X-0004609Y0005433D01*
Y0005520D01*
X-0004653Y0005608D01*
X-0004784D01*
X-0005007Y0005477D02*
X-0005138D01*
X-0004963Y0005345D02*
X-0005138D01*
Y0005608D01*
X-0004963D01*
X-0005317Y0005345D02*
X-0005470D01*
Y0005608D01*
X-0008861Y0004267D02*
X-0008839Y0004223D01*
X-0008708D01*
X-0008686Y0004267D01*
Y0004355D01*
X-0008730Y0004398D01*
X-0008861D01*
Y0004486D01*
X-0008686D01*
X-0009040Y0004223D02*
X-0009128D01*
X-0009084D02*
Y0004486D01*
X-0009128Y0004442D01*
X-0009350Y0004486D02*
Y0004267D01*
X-0009372Y0004223D01*
X-0009504D01*
X-0009526Y0004267D01*
Y0004486D01*
X0032678Y-0033174D02*
X0032546D01*
X0032524Y-0033130D01*
Y-0033086D01*
X0032546Y-0033042D01*
X0032678D01*
X0032700Y-0033086D01*
Y-0033130D01*
X0032612Y-0033305D01*
X0032988Y-0033042D02*
X0033032Y-0033086D01*
X0033054Y-0033130D01*
Y-0033217D01*
X0033032Y-0033261D01*
X0032988Y-0033305D01*
X0032944D01*
X0032901Y-0033261D01*
X0032879Y-0033217D01*
Y-0033130D01*
X0032901Y-0033086D01*
X0032944Y-0033042D01*
X0032988D01*
X0033233D02*
X0033320D01*
X0033277D02*
Y-0033305D01*
X0033320Y-0033261D01*
X0033543Y-0033305D02*
Y-0033217D01*
X0033631Y-0033042D01*
X0033719Y-0033217D01*
Y-0033305D01*
X0034073Y-0033174D02*
X0033942D01*
X0033898Y-0033217D01*
Y-0033261D01*
X0033942Y-0033305D01*
X0034073D01*
Y-0033042D01*
X-0016757Y0005477D02*
X-0016735Y0005520D01*
Y0005564D01*
X-0016757Y0005608D01*
X-0016888D01*
X-0016910Y0005564D01*
Y0005520D01*
X-0016888Y0005477D01*
X-0016757D01*
X-0016735Y0005433D01*
Y0005389D01*
X-0016757Y0005345D01*
X-0016888D01*
X-0016910Y0005389D01*
Y0005433D01*
X-0016888Y0005477D01*
X-0017089Y0005345D02*
X-0017264D01*
X-0017089Y0005520D01*
Y0005564D01*
X-0017111Y0005608D01*
X-0017242D01*
X-0017264Y0005564D01*
X-0017596Y0005345D02*
Y0005608D01*
X-0017619Y0005345D02*
X-0017487D01*
X-0017443Y0005433D01*
Y0005520D01*
X-0017487Y0005608D01*
X-0017619D01*
X-0017842Y0005477D02*
X-0017973D01*
X-0017798Y0005345D02*
X-0017973D01*
Y0005608D01*
X-0017798D01*
X-0018152Y0005345D02*
X-0018305D01*
Y0005608D01*
X0037156Y-0032657D02*
Y-0032482D01*
X0037331Y-0032657D01*
X0037375D01*
X0037419Y-0032635D01*
Y-0032504D01*
X0037375Y-0032482D01*
X0037419Y-0032303D02*
X0037331D01*
X0037156Y-0032215D01*
X0037331Y-0032128D01*
X0037419D01*
X0037288Y-0031774D02*
Y-0031905D01*
X0037331Y-0031949D01*
X0037375D01*
X0037419Y-0031905D01*
Y-0031774D01*
X0037156D01*
X0007027Y0005389D02*
X0007049Y0005345D01*
X0007180D01*
X0007202Y0005389D01*
Y0005477D01*
X0007158Y0005520D01*
X0007027D01*
Y0005608D01*
X0007202D01*
X0006848Y0005345D02*
X0006673D01*
X0006848Y0005520D01*
Y0005564D01*
X0006826Y0005608D01*
X0006695D01*
X0006673Y0005564D01*
X0006341Y0005345D02*
Y0005608D01*
X0006319Y0005345D02*
X0006450D01*
X0006494Y0005433D01*
Y0005520D01*
X0006450Y0005608D01*
X0006319D01*
X0006095Y0005477D02*
X0005964D01*
X0006139Y0005345D02*
X0005964D01*
Y0005608D01*
X0006139D01*
X0005785Y0005345D02*
X0005632D01*
Y0005608D01*
X0002241Y0004287D02*
X0002285Y0004243D01*
X0002372D01*
X0002417Y0004287D01*
Y0004331D01*
X0002329Y0004418D01*
X0002417Y0004506D01*
X0002241D01*
X0002062Y0004243D02*
X0001975D01*
X0002019D02*
Y0004506D01*
X0001975Y0004462D01*
X0001752Y0004506D02*
Y0004287D01*
X0001730Y0004243D01*
X0001599D01*
X0001577Y0004287D01*
Y0004506D01*
X-0008226Y-0033515D02*
X-0008139D01*
X-0007964Y-0033603D01*
X-0008139Y-0033690D01*
X-0008226D01*
X-0008007Y-0034044D02*
X-0007964Y-0034022D01*
Y-0033891D01*
X-0008007Y-0033869D01*
X-0008095D01*
X-0008139Y-0033913D01*
Y-0034044D01*
X-0008226D01*
Y-0033869D01*
X0034127Y-0032791D02*
X0034149Y-0032747D01*
Y-0032704D01*
X0034127Y-0032660D01*
X0033996D01*
X0033974Y-0032704D01*
Y-0032747D01*
X0033996Y-0032791D01*
X0034127D01*
X0034149Y-0032835D01*
Y-0032879D01*
X0034127Y-0032922D01*
X0033996D01*
X0033974Y-0032879D01*
Y-0032835D01*
X0033996Y-0032791D01*
X0033685Y-0032922D02*
X0033641Y-0032879D01*
X0033619Y-0032835D01*
Y-0032747D01*
X0033641Y-0032704D01*
X0033685Y-0032660D01*
X0033729D01*
X0033772Y-0032704D01*
X0033794Y-0032747D01*
Y-0032835D01*
X0033772Y-0032879D01*
X0033729Y-0032922D01*
X0033685D01*
X0033440D02*
X0033353D01*
X0033396D02*
Y-0032660D01*
X0033353Y-0032704D01*
X0033130Y-0032660D02*
Y-0032747D01*
X0033042Y-0032922D01*
X0032955Y-0032747D01*
Y-0032660D01*
X0032600Y-0032791D02*
X0032731D01*
X0032776Y-0032747D01*
Y-0032704D01*
X0032731Y-0032660D01*
X0032600D01*
Y-0032922D01*
X0016572Y0005413D02*
X0016397D01*
X0016485Y0005588D01*
X0016528D01*
Y0005326D01*
X0016218D02*
X0016043D01*
X0016218Y0005501D01*
Y0005544D01*
X0016196Y0005588D01*
X0016065D01*
X0016043Y0005544D01*
X0015711Y0005326D02*
Y0005588D01*
X0015689Y0005326D02*
X0015820D01*
X0015864Y0005413D01*
Y0005501D01*
X0015820Y0005588D01*
X0015689D01*
X0015465Y0005457D02*
X0015334D01*
X0015509Y0005326D02*
X0015334D01*
Y0005588D01*
X0015509D01*
X0015155Y0005326D02*
X0015002D01*
Y0005588D01*
X0018130Y0005369D02*
X0018173Y0005326D01*
X0018261D01*
X0018305Y0005369D01*
Y0005413D01*
X0018217Y0005501D01*
X0018305Y0005588D01*
X0018130D01*
X0017950Y0005326D02*
X0017775D01*
X0017950Y0005501D01*
Y0005544D01*
X0017928Y0005588D01*
X0017797D01*
X0017775Y0005544D01*
X0017443Y0005326D02*
Y0005588D01*
X0017421Y0005326D02*
X0017552D01*
X0017596Y0005413D01*
Y0005501D01*
X0017552Y0005588D01*
X0017421D01*
X0017198Y0005457D02*
X0017067D01*
X0017242Y0005326D02*
X0017067D01*
Y0005588D01*
X0017242D01*
X0016887Y0005326D02*
X0016734D01*
Y0005588D01*
X0013519Y0004243D02*
X0013344D01*
X0013519Y0004418D01*
Y0004462D01*
X0013497Y0004506D01*
X0013366D01*
X0013344Y0004462D01*
X0013165Y0004243D02*
X0013077D01*
X0013121D02*
Y0004506D01*
X0013077Y0004462D01*
X0012854Y0004506D02*
Y0004287D01*
X0012832Y0004243D01*
X0012701D01*
X0012679Y0004287D01*
Y0004506D01*
X0036008Y-0032517D02*
X0036052Y-0032539D01*
X0036096D01*
X0036139Y-0032517D01*
Y-0032386D01*
X0036096Y-0032364D01*
X0036052D01*
X0036008Y-0032386D01*
Y-0032517D01*
X0035965Y-0032539D01*
X0035920D01*
X0035877Y-0032517D01*
Y-0032386D01*
X0035920Y-0032364D01*
X0035965D01*
X0036008Y-0032386D01*
X0036139Y-0032185D02*
X0036052D01*
X0035877Y-0032097D01*
X0036052Y-0032010D01*
X0036139D01*
X0036008Y-0031656D02*
Y-0031787D01*
X0036052Y-0031831D01*
X0036096D01*
X0036139Y-0031787D01*
Y-0031656D01*
X0035877D01*
X0005317Y0005477D02*
X0005448D01*
X0005470Y0005433D01*
Y0005389D01*
X0005448Y0005345D01*
X0005317D01*
X0005295Y0005389D01*
Y0005433D01*
X0005382Y0005608D01*
X0005116Y0005345D02*
X0004941D01*
X0005116Y0005520D01*
Y0005564D01*
X0005094Y0005608D01*
X0004963D01*
X0004941Y0005564D01*
X0004608Y0005345D02*
Y0005608D01*
X0004586Y0005345D02*
X0004717D01*
X0004761Y0005433D01*
Y0005520D01*
X0004717Y0005608D01*
X0004586D01*
X0004363Y0005477D02*
X0004232D01*
X0004407Y0005345D02*
X0004232D01*
Y0005608D01*
X0004407D01*
X0004053Y0005345D02*
X0003900D01*
Y0005608D01*
X-0010354Y-0034730D02*
X-0010288Y-0034861D01*
X-0010463Y-0034730D02*
X-0010332D01*
X-0010288Y-0034686D01*
Y-0034643D01*
X-0010332Y-0034599D01*
X-0010463D01*
Y-0034861D01*
X-0010686Y-0034730D02*
X-0010817D01*
X-0010642Y-0034861D02*
X-0010817D01*
Y-0034599D01*
X-0010642D01*
X-0011150Y-0034861D02*
Y-0034599D01*
X-0011172Y-0034861D02*
X-0011041D01*
X-0010996Y-0034774D01*
Y-0034686D01*
X-0011041Y-0034599D01*
X-0011172D01*
X-0011351Y-0034774D02*
X-0011526D01*
X-0011351Y-0034861D02*
Y-0034730D01*
X-0011417Y-0034599D01*
X-0011460D01*
X-0011526Y-0034730D01*
Y-0034861D01*
X-0011749Y-0034730D02*
X-0011880D01*
X-0011705Y-0034861D02*
X-0011880D01*
Y-0034599D01*
X-0011705D01*
X-0012059Y-0034730D02*
X-0012235D01*
X-0012059Y-0034861D02*
Y-0034599D01*
X-0012235Y-0034861D02*
Y-0034599D01*
X-0013020Y-0034861D02*
Y-0034599D01*
X-0013042Y-0034861D02*
X-0012911D01*
X-0012867Y-0034774D01*
Y-0034686D01*
X-0012911Y-0034599D01*
X-0013042D01*
X-0013265Y-0034730D02*
X-0013396D01*
X-0013221Y-0034861D02*
X-0013396D01*
Y-0034599D01*
X-0013221D01*
X-0013575Y-0034861D02*
X-0013728D01*
Y-0034599D01*
X0013099Y0026428D02*
X0013056Y0026472D01*
X0013033Y0026516D01*
Y0026603D01*
X0013056Y0026647D01*
X0013099Y0026691D01*
X0013143D01*
X0013187Y0026647D01*
X0013209Y0026603D01*
Y0026516D01*
X0013187Y0026472D01*
X0013143Y0026428D01*
X0013099D01*
X0012854Y0026691D02*
Y0026472D01*
X0012832Y0026428D01*
X0012701D01*
X0012679Y0026472D01*
Y0026691D01*
X0007027Y-0005757D02*
X0007158Y-0005494D01*
X0006983D01*
X0006804Y-0005757D02*
X0006717D01*
X0006760D02*
Y-0005494D01*
X0006717Y-0005538D01*
X0006341Y-0005757D02*
Y-0005494D01*
X0006319Y-0005757D02*
X0006450D01*
X0006494Y-0005669D01*
Y-0005582D01*
X0006450Y-0005494D01*
X0006319D01*
X0006095Y-0005626D02*
X0005964D01*
X0006139Y-0005757D02*
X0005964D01*
Y-0005494D01*
X0006139D01*
X0005785Y-0005757D02*
X0005632D01*
Y-0005494D01*
X-0008928Y-0033314D02*
X-0009191D01*
X-0008928Y-0033336D02*
Y-0033205D01*
X-0009016Y-0033161D01*
X-0009104D01*
X-0009191Y-0033205D01*
Y-0033336D01*
Y-0033515D02*
X-0008928D01*
X-0008972Y-0033559D01*
X-0009147Y-0033646D01*
X-0009191Y-0033690D01*
X-0008928D01*
X-0009060Y-0033957D02*
Y-0033869D01*
X-0008972D01*
X-0008928Y-0033891D01*
Y-0034022D01*
X-0008972Y-0034044D01*
X-0009147D01*
X-0009191Y-0034022D01*
Y-0033891D01*
X-0009147Y-0033869D01*
X0002084Y-0006728D02*
X0001953D01*
X0001931Y-0006684D01*
Y-0006641D01*
X0001953Y-0006597D01*
X0002084D01*
X0002106Y-0006641D01*
Y-0006684D01*
X0002019Y-0006859D01*
X0001752Y-0006597D02*
Y-0006816D01*
X0001730Y-0006859D01*
X0001599D01*
X0001577Y-0006816D01*
Y-0006597D01*
X0034481Y-0032673D02*
X0034350D01*
X0034328Y-0032629D01*
Y-0032585D01*
X0034350Y-0032542D01*
X0034481D01*
X0034503Y-0032585D01*
Y-0032629D01*
X0034415Y-0032804D01*
X0034039D02*
X0033996Y-0032761D01*
X0033974Y-0032717D01*
Y-0032629D01*
X0033996Y-0032585D01*
X0034039Y-0032542D01*
X0034083D01*
X0034127Y-0032585D01*
X0034149Y-0032629D01*
Y-0032717D01*
X0034127Y-0032761D01*
X0034083Y-0032804D01*
X0034039D01*
X0033794D02*
X0033707D01*
X0033751D02*
Y-0032542D01*
X0033707Y-0032585D01*
X0033484Y-0032542D02*
Y-0032629D01*
X0033396Y-0032804D01*
X0033309Y-0032629D01*
Y-0032542D01*
X0032955Y-0032673D02*
X0033086D01*
X0033130Y-0032629D01*
Y-0032585D01*
X0033086Y-0032542D01*
X0032955D01*
Y-0032804D01*
X0036664Y-0032889D02*
Y-0032802D01*
Y-0032845D02*
X0036927D01*
X0036883Y-0032802D01*
X0036927Y-0032579D02*
X0036839D01*
X0036664Y-0032491D01*
X0036839Y-0032404D01*
X0036927D01*
X0036796Y-0032049D02*
Y-0032180D01*
X0036839Y-0032224D01*
X0036883D01*
X0036927Y-0032180D01*
Y-0032049D01*
X0036664D01*
X-0016844Y-0005757D02*
X-0016888Y-0005713D01*
X-0016910Y-0005669D01*
Y-0005582D01*
X-0016888Y-0005538D01*
X-0016844Y-0005494D01*
X-0016800D01*
X-0016757Y-0005538D01*
X-0016735Y-0005582D01*
Y-0005669D01*
X-0016757Y-0005713D01*
X-0016800Y-0005757D01*
X-0016844D01*
X-0017089D02*
X-0017264D01*
X-0017089Y-0005582D01*
Y-0005538D01*
X-0017111Y-0005494D01*
X-0017242D01*
X-0017264Y-0005538D01*
X-0017596Y-0005757D02*
Y-0005494D01*
X-0017619Y-0005757D02*
X-0017487D01*
X-0017443Y-0005669D01*
Y-0005582D01*
X-0017487Y-0005494D01*
X-0017619D01*
X-0017842Y-0005626D02*
X-0017973D01*
X-0017798Y-0005757D02*
X-0017973D01*
Y-0005494D01*
X-0017798D01*
X-0018152Y-0005757D02*
X-0018305D01*
Y-0005494D01*
X-0015049Y-0005626D02*
X-0015180D01*
X-0015202Y-0005582D01*
Y-0005538D01*
X-0015180Y-0005494D01*
X-0015049D01*
X-0015027Y-0005538D01*
Y-0005582D01*
X-0015115Y-0005757D01*
X-0015381D02*
X-0015469D01*
X-0015425D02*
Y-0005494D01*
X-0015469Y-0005538D01*
X-0015844Y-0005757D02*
Y-0005494D01*
X-0015867Y-0005757D02*
X-0015735D01*
X-0015691Y-0005669D01*
Y-0005582D01*
X-0015735Y-0005494D01*
X-0015867D01*
X-0016090Y-0005626D02*
X-0016221D01*
X-0016046Y-0005757D02*
X-0016221D01*
Y-0005494D01*
X-0016046D01*
X-0016400Y-0005757D02*
X-0016553D01*
Y-0005494D01*
X0034589Y-0032771D02*
X0034546Y-0032727D01*
X0034458D01*
X0034414Y-0032771D01*
Y-0032815D01*
X0034502Y-0032902D01*
X0034414Y-0032990D01*
X0034589D01*
X0034878Y-0032727D02*
X0034922Y-0032771D01*
X0034944Y-0032815D01*
Y-0032902D01*
X0034922Y-0032946D01*
X0034878Y-0032990D01*
X0034834D01*
X0034791Y-0032946D01*
X0034769Y-0032902D01*
Y-0032815D01*
X0034791Y-0032771D01*
X0034834Y-0032727D01*
X0034878D01*
X0035123D02*
X0035210D01*
X0035167D02*
Y-0032990D01*
X0035210Y-0032946D01*
X0035433Y-0032990D02*
Y-0032902D01*
X0035521Y-0032727D01*
X0035608Y-0032902D01*
Y-0032990D01*
X0035963Y-0032859D02*
X0035831D01*
X0035787Y-0032902D01*
Y-0032946D01*
X0035831Y-0032990D01*
X0035963D01*
Y-0032727D01*
X0037333Y-0034241D02*
X0037246D01*
X0037289D02*
Y-0033979D01*
X0037246Y-0034022D01*
X0037023Y-0034241D02*
X0036848D01*
X0037023Y-0034066D01*
Y-0034022D01*
X0037001Y-0033979D01*
X0036870D01*
X0036848Y-0034022D01*
X0036669Y-0034241D02*
X0036581D01*
X0036625D02*
Y-0033979D01*
X0036581Y-0034022D01*
X0036358Y-0033979D02*
Y-0034066D01*
X0036270Y-0034241D01*
X0036183Y-0034066D01*
Y-0033979D01*
X0035829Y-0034110D02*
X0035960D01*
X0036004Y-0034066D01*
Y-0034022D01*
X0035960Y-0033979D01*
X0035829D01*
Y-0034241D01*
X0038291Y-0032194D02*
X0038248Y-0032150D01*
X0038226Y-0032106D01*
Y-0032019D01*
X0038248Y-0031975D01*
X0038291Y-0031931D01*
X0038335D01*
X0038379Y-0031975D01*
X0038401Y-0032019D01*
Y-0032106D01*
X0038379Y-0032150D01*
X0038335Y-0032194D01*
X0038291D01*
X0038046D02*
X0037871D01*
X0038046Y-0032019D01*
Y-0031975D01*
X0038024Y-0031931D01*
X0037893D01*
X0037871Y-0031975D01*
X0037692Y-0032194D02*
X0037605D01*
X0037648D02*
Y-0031931D01*
X0037605Y-0031975D01*
X0037382Y-0031931D02*
Y-0032019D01*
X0037294Y-0032194D01*
X0037207Y-0032019D01*
Y-0031931D01*
X0036852Y-0032063D02*
X0036983D01*
X0037028Y-0032019D01*
Y-0031975D01*
X0036983Y-0031931D01*
X0036852D01*
Y-0032194D01*
X-0019898Y-0006859D02*
X-0019941Y-0006816D01*
X-0019963Y-0006772D01*
Y-0006684D01*
X-0019941Y-0006641D01*
X-0019898Y-0006597D01*
X-0019854D01*
X-0019810Y-0006641D01*
X-0019788Y-0006684D01*
Y-0006772D01*
X-0019810Y-0006816D01*
X-0019854Y-0006859D01*
X-0019898D01*
X-0020143D02*
X-0020230D01*
X-0020186D02*
Y-0006597D01*
X-0020230Y-0006641D01*
X-0020453Y-0006597D02*
Y-0006816D01*
X-0020475Y-0006859D01*
X-0020606D01*
X-0020628Y-0006816D01*
Y-0006597D01*
X-0005632Y-0005757D02*
X-0005807D01*
X-0005632Y-0005582D01*
Y-0005538D01*
X-0005654Y-0005494D01*
X-0005785D01*
X-0005807Y-0005538D01*
X-0005987Y-0005757D02*
X-0006162D01*
X-0005987Y-0005582D01*
Y-0005538D01*
X-0006009Y-0005494D01*
X-0006140D01*
X-0006162Y-0005538D01*
X-0006494Y-0005757D02*
Y-0005494D01*
X-0006516Y-0005757D02*
X-0006385D01*
X-0006341Y-0005669D01*
Y-0005582D01*
X-0006385Y-0005494D01*
X-0006516D01*
X-0006739Y-0005626D02*
X-0006870D01*
X-0006695Y-0005757D02*
X-0006870D01*
Y-0005494D01*
X-0006695D01*
X-0007050Y-0005757D02*
X-0007203D01*
Y-0005494D01*
X0036799Y-0034110D02*
X0036668D01*
X0036646Y-0034066D01*
Y-0034022D01*
X0036668Y-0033979D01*
X0036799D01*
X0036821Y-0034022D01*
Y-0034066D01*
X0036733Y-0034241D01*
X0036467D02*
X0036380D01*
X0036423D02*
Y-0033979D01*
X0036380Y-0034022D01*
X0036157Y-0034241D02*
X0036069D01*
X0036113D02*
Y-0033979D01*
X0036069Y-0034022D01*
X0035846Y-0033979D02*
Y-0034066D01*
X0035759Y-0034241D01*
X0035671Y-0034066D01*
Y-0033979D01*
X0035317Y-0034110D02*
X0035448D01*
X0035492Y-0034066D01*
Y-0034022D01*
X0035448Y-0033979D01*
X0035317D01*
Y-0034241D01*
X0034665Y-0030656D02*
X0034507D01*
X0034481Y-0030604D01*
Y-0030551D01*
X0034507Y-0030499D01*
X0034665D01*
X0034691Y-0030551D01*
Y-0030604D01*
X0034586Y-0030814D01*
X0034087Y-0030761D02*
X0034114Y-0030814D01*
X0034271D01*
X0034298Y-0030761D01*
Y-0030656D01*
X0034245Y-0030604D01*
X0034087D01*
Y-0030499D01*
X0034298D01*
X0033904Y-0030814D02*
X0033799D01*
X0033852D02*
Y-0030499D01*
X0033799Y-0030551D01*
X0033563Y-0030499D02*
Y-0030604D01*
X0033458Y-0030814D01*
X0033353Y-0030604D01*
Y-0030499D01*
X0032959Y-0030656D02*
X0033117D01*
X0033169Y-0030604D01*
Y-0030551D01*
X0033117Y-0030499D01*
X0032959D01*
Y-0030814D01*
X0034626Y-0031148D02*
X0034652Y-0031096D01*
Y-0031043D01*
X0034626Y-0030991D01*
X0034468D01*
X0034442Y-0031043D01*
Y-0031096D01*
X0034468Y-0031148D01*
X0034626D01*
X0034652Y-0031201D01*
Y-0031254D01*
X0034626Y-0031306D01*
X0034468D01*
X0034442Y-0031254D01*
Y-0031201D01*
X0034468Y-0031148D01*
X0034048Y-0031254D02*
X0034074Y-0031306D01*
X0034232D01*
X0034258Y-0031254D01*
Y-0031148D01*
X0034206Y-0031096D01*
X0034048D01*
Y-0030991D01*
X0034258D01*
X0033865Y-0031306D02*
X0033760D01*
X0033812D02*
Y-0030991D01*
X0033760Y-0031043D01*
X0033524Y-0030991D02*
Y-0031096D01*
X0033419Y-0031306D01*
X0033313Y-0031096D01*
Y-0030991D01*
X0032920Y-0031148D02*
X0033077D01*
X0033130Y-0031096D01*
Y-0031043D01*
X0033077Y-0030991D01*
X0032920D01*
Y-0031306D01*
X0032856Y-0031407D02*
X0032987Y-0031144D01*
X0032812D01*
X0032633Y-0031319D02*
X0032458D01*
X0032545Y-0031144D01*
X0032589D01*
Y-0031407D01*
X0032279D02*
X0032191D01*
X0032235D02*
Y-0031144D01*
X0032191Y-0031188D01*
X0031969Y-0031144D02*
Y-0031231D01*
X0031881Y-0031407D01*
X0031793Y-0031231D01*
Y-0031144D01*
X0031439Y-0031275D02*
X0031570D01*
X0031614Y-0031231D01*
Y-0031188D01*
X0031570Y-0031144D01*
X0031439D01*
Y-0031407D01*
X0034737Y-0031748D02*
X0034759Y-0031704D01*
Y-0031660D01*
X0034737Y-0031617D01*
X0034606D01*
X0034584Y-0031660D01*
Y-0031704D01*
X0034606Y-0031748D01*
X0034737D01*
X0034759Y-0031791D01*
Y-0031835D01*
X0034737Y-0031879D01*
X0034606D01*
X0034584Y-0031835D01*
Y-0031791D01*
X0034606Y-0031748D01*
X0034405Y-0031791D02*
X0034230D01*
X0034317Y-0031617D01*
X0034361D01*
Y-0031879D01*
X0034050D02*
X0033963D01*
X0034007D02*
Y-0031617D01*
X0033963Y-0031660D01*
X0033740Y-0031617D02*
Y-0031704D01*
X0033652Y-0031879D01*
X0033565Y-0031704D01*
Y-0031617D01*
X0033211Y-0031748D02*
X0033342D01*
X0033386Y-0031704D01*
Y-0031660D01*
X0033342Y-0031617D01*
X0033211D01*
Y-0031879D01*
X0056003Y0035120D02*
X0056090Y0035295D01*
Y0035470D01*
X0056003Y0035645D01*
X0055408Y0035120D02*
Y0035645D01*
X0055364Y0035120D02*
X0055626D01*
X0055714Y0035295D01*
Y0035470D01*
X0055626Y0035645D01*
X0055364D01*
X0055163Y0035295D02*
X0054813D01*
X0055163Y0035120D02*
Y0035383D01*
X0055031Y0035645D01*
X0054944D01*
X0054813Y0035383D01*
Y0035120D01*
X0054262Y0035383D02*
X0054524D01*
X0054612Y0035470D01*
Y0035557D01*
X0054524Y0035645D01*
X0054262D01*
Y0035120D01*
X0054061D02*
X0053886D01*
X0053973D02*
Y0035645D01*
X0054061D02*
X0053886D01*
X0053422Y0035120D02*
Y0035645D01*
X0053597D02*
X0053247D01*
X0053046D02*
Y0035120D01*
X0052958Y0035207D01*
X0052783Y0035557D01*
X0052696Y0035645D01*
Y0035120D01*
X0052495Y0035295D02*
X0052145D01*
X0052495Y0035120D02*
Y0035383D01*
X0052363Y0035645D01*
X0052276D01*
X0052145Y0035383D01*
Y0035120D01*
X0051108Y0035383D02*
X0050846D01*
X0051196Y0035120D02*
X0050846D01*
Y0035645D01*
X0051196D01*
X0050644D02*
Y0035120D01*
X0050557Y0035207D01*
X0050382Y0035557D01*
X0050294Y0035645D01*
Y0035120D01*
X0050093Y0035295D02*
X0049743D01*
X0050093Y0035120D02*
Y0035383D01*
X0049962Y0035645D01*
X0049874D01*
X0049743Y0035383D01*
Y0035120D01*
X0049542D02*
X0049236D01*
Y0035645D01*
X0048685Y0035383D02*
X0048947D01*
X0049035Y0035470D01*
Y0035557D01*
X0048947Y0035645D01*
X0048685D01*
Y0035120D01*
X0047736D02*
Y0035645D01*
X0047648Y0035557D01*
X0047561Y0035383D01*
X0047473Y0035557D01*
X0047386Y0035645D01*
Y0035120D01*
X0047185D02*
Y0035645D01*
X0047097Y0035557D01*
X0047009Y0035383D01*
X0046922Y0035557D01*
X0046835Y0035645D01*
Y0035120D01*
X0046283Y0035207D02*
X0046327Y0035120D01*
X0046589D01*
X0046633Y0035207D01*
Y0035383D01*
X0046546Y0035470D01*
X0046283D01*
Y0035645D01*
X0046633D01*
X0045732Y0035207D02*
X0045776Y0035120D01*
X0046038D01*
X0046082Y0035207D01*
Y0035383D01*
X0045994Y0035470D01*
X0045732D01*
Y0035645D01*
X0046082D01*
X0045444Y0035120D02*
X0045531D01*
Y0035207D01*
X0045444D01*
Y0035120D01*
X0044936D02*
X0044849Y0035207D01*
X0044805Y0035295D01*
Y0035470D01*
X0044849Y0035557D01*
X0044936Y0035645D01*
X0045024D01*
X0045111Y0035557D01*
X0045155Y0035470D01*
Y0035295D01*
X0045111Y0035207D01*
X0045024Y0035120D01*
X0044936D01*
X0044604D02*
X0044517Y0035295D01*
Y0035470D01*
X0044604Y0035645D01*
X0043305Y0035383D02*
X0043043D01*
X0043393Y0035120D02*
X0043043D01*
Y0035645D01*
X0043393D01*
X0042841Y0035120D02*
X0042535D01*
Y0035645D01*
X0042028Y0035120D02*
X0041984Y0035207D01*
Y0035557D01*
X0042028Y0035645D01*
X0042290D01*
X0042334Y0035557D01*
Y0035207D01*
X0042290Y0035120D01*
X0042028D01*
X0041783Y0035383D02*
X0041433D01*
X0041783Y0035120D02*
Y0035645D01*
X0041433Y0035120D02*
Y0035645D01*
X0040484Y0035120D02*
Y0035645D01*
X0040396Y0035557D01*
X0040309Y0035383D01*
X0040221Y0035557D01*
X0040134Y0035645D01*
Y0035120D01*
X0039933D02*
Y0035645D01*
X0039845Y0035557D01*
X0039757Y0035383D01*
X0039670Y0035557D01*
X0039583Y0035645D01*
Y0035120D01*
X0039031Y0035207D02*
X0039075Y0035120D01*
X0039337D01*
X0039381Y0035207D01*
Y0035383D01*
X0039294Y0035470D01*
X0039031D01*
Y0035645D01*
X0039381D01*
X0038830Y0035120D02*
X0038656D01*
X0038743D02*
Y0035645D01*
X0038656Y0035557D01*
X0038280Y0035120D02*
X0038367D01*
Y0035207D01*
X0038280D01*
Y0035120D01*
X0037772D02*
X0037685Y0035207D01*
X0037641Y0035295D01*
Y0035470D01*
X0037685Y0035557D01*
X0037772Y0035645D01*
X0037859D01*
X0037947Y0035557D01*
X0037991Y0035470D01*
Y0035295D01*
X0037947Y0035207D01*
X0037859Y0035120D01*
X0037772D01*
X0036692Y0035645D02*
X0036430Y0035120D01*
X0035130D02*
Y0035645D01*
X0035087Y0035120D02*
X0035349D01*
X0035437Y0035295D01*
Y0035470D01*
X0035349Y0035645D01*
X0035087D01*
X0034885Y0035295D02*
X0034535D01*
X0034885Y0035120D02*
Y0035383D01*
X0034754Y0035645D01*
X0034667D01*
X0034535Y0035383D01*
Y0035120D01*
X0033984Y0035383D02*
X0034246D01*
X0034334Y0035470D01*
Y0035557D01*
X0034246Y0035645D01*
X0033984D01*
Y0035120D01*
X0033035D02*
Y0035645D01*
X0032947Y0035557D01*
X0032860Y0035383D01*
X0032772Y0035557D01*
X0032685Y0035645D01*
Y0035120D01*
X0032484D02*
Y0035645D01*
X0032396Y0035557D01*
X0032309Y0035383D01*
X0032221Y0035557D01*
X0032134Y0035645D01*
Y0035120D01*
X0031933Y0035295D02*
X0031583D01*
X0031757Y0035645D01*
X0031845D01*
Y0035120D01*
X0031294D02*
X0031381D01*
Y0035207D01*
X0031294D01*
Y0035120D01*
X0030787D02*
X0030699Y0035207D01*
X0030656Y0035295D01*
Y0035470D01*
X0030699Y0035557D01*
X0030787Y0035645D01*
X0030874D01*
X0030961Y0035557D01*
X0031006Y0035470D01*
Y0035295D01*
X0030961Y0035207D01*
X0030874Y0035120D01*
X0030787D01*
X0029706Y0035383D02*
X0029356D01*
X0028407Y0035120D02*
X0028232D01*
X0028320D02*
Y0035645D01*
X0028232Y0035557D01*
X0027944Y0035295D02*
X0027594D01*
X0027944Y0035120D02*
Y0035383D01*
X0027812Y0035645D01*
X0027725D01*
X0027594Y0035383D01*
Y0035120D01*
X0027393D02*
X0027218D01*
X0027305D02*
Y0035645D01*
X0027393D02*
X0027218D01*
X0026929D02*
Y0035470D01*
X0026754Y0035120D01*
X0026579Y0035470D01*
Y0035645D01*
X-0003944Y-0005757D02*
X-0004031D01*
X-0003988D02*
Y-0005494D01*
X-0004031Y-0005538D01*
X-0004254Y-0005757D02*
X-0004430D01*
X-0004254Y-0005582D01*
Y-0005538D01*
X-0004276Y-0005494D01*
X-0004407D01*
X-0004430Y-0005538D01*
X-0004762Y-0005757D02*
Y-0005494D01*
X-0004784Y-0005757D02*
X-0004653D01*
X-0004609Y-0005669D01*
Y-0005582D01*
X-0004653Y-0005494D01*
X-0004784D01*
X-0005007Y-0005626D02*
X-0005138D01*
X-0004963Y-0005757D02*
X-0005138D01*
Y-0005494D01*
X-0004963D01*
X-0005317Y-0005757D02*
X-0005470D01*
Y-0005494D01*
X0016572Y0027638D02*
X0016397D01*
X0016485Y0027813D01*
X0016528D01*
Y0027550D01*
X0016043Y0027594D02*
X0016087Y0027550D01*
X0016174D01*
X0016218Y0027594D01*
Y0027638D01*
X0016130Y0027725D01*
X0016218Y0027813D01*
X0016043D01*
X0015711Y0027550D02*
Y0027813D01*
X0015689Y0027550D02*
X0015820D01*
X0015864Y0027638D01*
Y0027725D01*
X0015820Y0027813D01*
X0015689D01*
X0015465Y0027681D02*
X0015334D01*
X0015509Y0027550D02*
X0015334D01*
Y0027813D01*
X0015509D01*
X0015155Y0027550D02*
X0015002D01*
Y0027813D01*
X-0008730Y-0006859D02*
X-0008817D01*
X-0008774D02*
Y-0006597D01*
X-0008817Y-0006641D01*
X-0009040Y-0006859D02*
X-0009128D01*
X-0009084D02*
Y-0006597D01*
X-0009128Y-0006641D01*
X-0009350Y-0006597D02*
Y-0006816D01*
X-0009372Y-0006859D01*
X-0009504D01*
X-0009526Y-0006816D01*
Y-0006597D01*
X0016415Y-0005606D02*
X0016546D01*
X0016568Y-0005650D01*
Y-0005694D01*
X0016546Y-0005737D01*
X0016415D01*
X0016393Y-0005694D01*
Y-0005650D01*
X0016480Y-0005475D01*
X0016213Y-0005737D02*
X0016126D01*
X0016170D02*
Y-0005475D01*
X0016126Y-0005519D01*
X0015750Y-0005737D02*
Y-0005475D01*
X0015728Y-0005737D02*
X0015859D01*
X0015903Y-0005650D01*
Y-0005562D01*
X0015859Y-0005475D01*
X0015728D01*
X0015505Y-0005606D02*
X0015374D01*
X0015549Y-0005737D02*
X0015374D01*
Y-0005475D01*
X0015549D01*
X0015194Y-0005737D02*
X0015041D01*
Y-0005475D01*
X0034997Y-0032957D02*
X0035041Y-0033001D01*
X0035128D01*
X0035172Y-0032957D01*
Y-0032913D01*
X0035085Y-0032826D01*
X0035172Y-0032739D01*
X0034997D01*
X0034643Y-0032957D02*
X0034665Y-0033001D01*
X0034796D01*
X0034818Y-0032957D01*
Y-0032870D01*
X0034774Y-0032826D01*
X0034643D01*
Y-0032739D01*
X0034818D01*
X0034464Y-0033001D02*
X0034376D01*
X0034420D02*
Y-0032739D01*
X0034376Y-0032782D01*
X0034154Y-0032739D02*
Y-0032826D01*
X0034066Y-0033001D01*
X0033978Y-0032826D01*
Y-0032739D01*
X0033624Y-0032870D02*
X0033755D01*
X0033799Y-0032826D01*
Y-0032782D01*
X0033755Y-0032739D01*
X0033624D01*
Y-0033001D01*
X0032594Y-0032174D02*
X0032419D01*
X0032594Y-0031999D01*
Y-0031956D01*
X0032572Y-0031912D01*
X0032441D01*
X0032419Y-0031956D01*
X0032239Y-0032087D02*
X0032064D01*
X0032152Y-0031912D01*
X0032195D01*
Y-0032174D01*
X0031885D02*
X0031798D01*
X0031841D02*
Y-0031912D01*
X0031798Y-0031956D01*
X0031575Y-0031912D02*
Y-0031999D01*
X0031487Y-0032174D01*
X0031400Y-0031999D01*
Y-0031912D01*
X0031045Y-0032043D02*
X0031176D01*
X0031220Y-0031999D01*
Y-0031956D01*
X0031176Y-0031912D01*
X0031045D01*
Y-0032174D01*
X0018085Y-0005694D02*
X0018107Y-0005737D01*
X0018239D01*
X0018261Y-0005694D01*
Y-0005606D01*
X0018217Y-0005562D01*
X0018085D01*
Y-0005475D01*
X0018261D01*
X0017906Y-0005737D02*
X0017819D01*
X0017863D02*
Y-0005475D01*
X0017819Y-0005519D01*
X0017443Y-0005737D02*
Y-0005475D01*
X0017421Y-0005737D02*
X0017552D01*
X0017596Y-0005650D01*
Y-0005562D01*
X0017552Y-0005475D01*
X0017421D01*
X0017198Y-0005606D02*
X0017067D01*
X0017242Y-0005737D02*
X0017067D01*
Y-0005475D01*
X0017242D01*
X0016887Y-0005737D02*
X0016734D01*
Y-0005475D01*
X0013187Y-0006748D02*
X0013209Y-0006704D01*
Y-0006660D01*
X0013187Y-0006617D01*
X0013056D01*
X0013033Y-0006660D01*
Y-0006704D01*
X0013056Y-0006748D01*
X0013187D01*
X0013209Y-0006791D01*
Y-0006835D01*
X0013187Y-0006879D01*
X0013056D01*
X0013033Y-0006835D01*
Y-0006791D01*
X0013056Y-0006748D01*
X0012854Y-0006617D02*
Y-0006835D01*
X0012832Y-0006879D01*
X0012701D01*
X0012679Y-0006835D01*
Y-0006617D01*
X0033005Y-0031708D02*
X0032874D01*
X0032852Y-0031665D01*
Y-0031621D01*
X0032874Y-0031577D01*
X0033005D01*
X0033027Y-0031621D01*
Y-0031665D01*
X0032939Y-0031840D01*
X0032672Y-0031752D02*
X0032497D01*
X0032585Y-0031577D01*
X0032628D01*
Y-0031840D01*
X0032318D02*
X0032231D01*
X0032274D02*
Y-0031577D01*
X0032231Y-0031621D01*
X0032008Y-0031577D02*
Y-0031665D01*
X0031920Y-0031840D01*
X0031833Y-0031665D01*
Y-0031577D01*
X0031478Y-0031708D02*
X0031609D01*
X0031654Y-0031665D01*
Y-0031621D01*
X0031609Y-0031577D01*
X0031478D01*
Y-0031840D01*
X0034645Y-0031236D02*
X0034776D01*
X0034798Y-0031280D01*
Y-0031324D01*
X0034776Y-0031367D01*
X0034645D01*
X0034623Y-0031324D01*
Y-0031280D01*
X0034711Y-0031105D01*
X0034444Y-0031280D02*
X0034269D01*
X0034356Y-0031105D01*
X0034400D01*
Y-0031367D01*
X0034090D02*
X0034002D01*
X0034046D02*
Y-0031105D01*
X0034002Y-0031148D01*
X0033780Y-0031105D02*
Y-0031192D01*
X0033692Y-0031367D01*
X0033604Y-0031192D01*
Y-0031105D01*
X0033250Y-0031236D02*
X0033381D01*
X0033425Y-0031192D01*
Y-0031148D01*
X0033381Y-0031105D01*
X0033250D01*
Y-0031367D01*
X0033115Y-0032224D02*
X0033290D01*
X0033203Y-0032399D01*
X0033159D01*
Y-0032137D01*
X0033579D02*
X0033622Y-0032180D01*
X0033644Y-0032224D01*
Y-0032312D01*
X0033622Y-0032356D01*
X0033579Y-0032399D01*
X0033535D01*
X0033491Y-0032356D01*
X0033469Y-0032312D01*
Y-0032224D01*
X0033491Y-0032180D01*
X0033535Y-0032137D01*
X0033579D01*
X0033824D02*
X0033911D01*
X0033867D02*
Y-0032399D01*
X0033911Y-0032356D01*
X0034134Y-0032399D02*
Y-0032312D01*
X0034222Y-0032137D01*
X0034309Y-0032312D01*
Y-0032399D01*
X0034663Y-0032268D02*
X0034532D01*
X0034488Y-0032312D01*
Y-0032356D01*
X0034532Y-0032399D01*
X0034663D01*
Y-0032137D01*
X0005443Y-0005626D02*
X0005465Y-0005582D01*
Y-0005538D01*
X0005443Y-0005494D01*
X0005312D01*
X0005290Y-0005538D01*
Y-0005582D01*
X0005312Y-0005626D01*
X0005443D01*
X0005465Y-0005669D01*
Y-0005713D01*
X0005443Y-0005757D01*
X0005312D01*
X0005290Y-0005713D01*
Y-0005669D01*
X0005312Y-0005626D01*
X0005111Y-0005757D02*
X0005024D01*
X0005067D02*
Y-0005494D01*
X0005024Y-0005538D01*
X0004648Y-0005757D02*
Y-0005494D01*
X0004626Y-0005757D02*
X0004757D01*
X0004801Y-0005669D01*
Y-0005582D01*
X0004757Y-0005494D01*
X0004626D01*
X0004402Y-0005626D02*
X0004271D01*
X0004446Y-0005757D02*
X0004271D01*
Y-0005494D01*
X0004446D01*
X0004092Y-0005757D02*
X0003939D01*
Y-0005494D01*
X0034317Y-0032881D02*
X0034213D01*
X0034265D02*
Y-0032566D01*
X0034213Y-0032618D01*
X0033976Y-0032723D02*
X0033766D01*
X0033976Y-0032881D02*
Y-0032566D01*
X0033766Y-0032881D02*
Y-0032566D01*
X0033478Y-0032881D02*
Y-0032566D01*
X0033583D02*
X0033372D01*
X0033189Y-0032881D02*
Y-0032566D01*
X0033136Y-0032618D01*
X0033084Y-0032723D01*
X0033031Y-0032618D01*
X0032979Y-0032566D01*
Y-0032881D01*
X0032795Y-0032828D02*
X0032769Y-0032881D01*
X0032611D01*
X0032585Y-0032828D01*
Y-0032618D01*
X0032611Y-0032566D01*
X0032769D01*
X0032795Y-0032618D01*
X0034587Y-0033137D02*
X0034376D01*
X0034587Y-0032927D01*
Y-0032874D01*
X0034560Y-0032822D01*
X0034403D01*
X0034376Y-0032874D01*
X0034193Y-0032979D02*
X0033983D01*
X0034193Y-0033137D02*
Y-0032822D01*
X0033983Y-0033137D02*
Y-0032822D01*
X0033694Y-0033137D02*
Y-0032822D01*
X0033799D02*
X0033589D01*
X0033406Y-0033137D02*
Y-0032822D01*
X0033353Y-0032874D01*
X0033300Y-0032979D01*
X0033248Y-0032874D01*
X0033195Y-0032822D01*
Y-0033137D01*
X0033012Y-0033084D02*
X0032985Y-0033137D01*
X0032828D01*
X0032802Y-0033084D01*
Y-0032874D01*
X0032828Y-0032822D01*
X0032985D01*
X0033012Y-0032874D01*
X-0015091Y0016448D02*
X-0015178D01*
X-0015134D02*
Y0016710D01*
X-0015178Y0016667D01*
X-0015401Y0016448D02*
X-0015488D01*
X-0015444D02*
Y0016710D01*
X-0015488Y0016667D01*
X-0015864Y0016448D02*
Y0016710D01*
X-0015886Y0016448D02*
X-0015755D01*
X-0015711Y0016535D01*
Y0016623D01*
X-0015755Y0016710D01*
X-0015886D01*
X-0016109Y0016579D02*
X-0016241D01*
X-0016065Y0016448D02*
X-0016241D01*
Y0016710D01*
X-0016065D01*
X-0016420Y0016448D02*
X-0016573D01*
Y0016710D01*
X0035437Y-0033375D02*
X0035393Y-0033331D01*
X0035371Y-0033287D01*
Y-0033200D01*
X0035393Y-0033156D01*
X0035437Y-0033113D01*
X0035481D01*
X0035524Y-0033156D01*
X0035546Y-0033200D01*
Y-0033287D01*
X0035524Y-0033331D01*
X0035481Y-0033375D01*
X0035437D01*
X0035017Y-0033331D02*
X0035039Y-0033375D01*
X0035170D01*
X0035192Y-0033331D01*
Y-0033244D01*
X0035148Y-0033200D01*
X0035017D01*
Y-0033113D01*
X0035192D01*
X0034838Y-0033375D02*
X0034750D01*
X0034794D02*
Y-0033113D01*
X0034750Y-0033156D01*
X0034528Y-0033113D02*
Y-0033200D01*
X0034440Y-0033375D01*
X0034352Y-0033200D01*
Y-0033113D01*
X0033998Y-0033244D02*
X0034129D01*
X0034173Y-0033200D01*
Y-0033156D01*
X0034129Y-0033113D01*
X0033998D01*
Y-0033375D01*
X0035128D02*
X0035041D01*
X0035085D02*
Y-0033113D01*
X0035041Y-0033156D01*
X0034643Y-0033331D02*
X0034665Y-0033375D01*
X0034796D01*
X0034818Y-0033331D01*
Y-0033244D01*
X0034774Y-0033200D01*
X0034643D01*
Y-0033113D01*
X0034818D01*
X0034464Y-0033375D02*
X0034376D01*
X0034420D02*
Y-0033113D01*
X0034376Y-0033156D01*
X0034154Y-0033113D02*
Y-0033200D01*
X0034066Y-0033375D01*
X0033978Y-0033200D01*
Y-0033113D01*
X0033624Y-0033244D02*
X0033755D01*
X0033799Y-0033200D01*
Y-0033156D01*
X0033755Y-0033113D01*
X0033624D01*
Y-0033375D01*
X-0020252Y0015457D02*
X-0020120D01*
X-0020098Y0015413D01*
Y0015369D01*
X-0020120Y0015326D01*
X-0020252D01*
X-0020274Y0015369D01*
Y0015413D01*
X-0020186Y0015588D01*
X-0020453D02*
Y0015369D01*
X-0020475Y0015326D01*
X-0020606D01*
X-0020628Y0015369D01*
Y0015588D01*
X0064479Y0022786D02*
Y0023049D01*
X0064567D02*
X0064392D01*
X0064213Y0023005D02*
X0064191Y0023049D01*
X0064059D01*
X0064037Y0023005D01*
Y0022961D01*
X0064059Y0022918D01*
X0064191D01*
X0064213Y0022874D01*
Y0022830D01*
X0064191Y0022786D01*
X0064059D01*
X0064037Y0022830D01*
X0063858Y0023005D02*
X0063836Y0023049D01*
X0063705D01*
X0063683Y0023005D01*
Y0022961D01*
X0063705Y0022918D01*
X0063836D01*
X0063858Y0022874D01*
Y0022830D01*
X0063836Y0022786D01*
X0063705D01*
X0063683Y0022830D01*
X-0005637Y0016535D02*
X-0005812D01*
X-0005725Y0016710D01*
X-0005681D01*
Y0016448D01*
X-0005991D02*
X-0006079D01*
X-0006035D02*
Y0016710D01*
X-0006079Y0016667D01*
X-0006455Y0016448D02*
Y0016710D01*
X-0006477Y0016448D02*
X-0006346D01*
X-0006302Y0016535D01*
Y0016623D01*
X-0006346Y0016710D01*
X-0006477D01*
X-0006700Y0016579D02*
X-0006831D01*
X-0006656Y0016448D02*
X-0006831D01*
Y0016710D01*
X-0006656D01*
X-0007010Y0016448D02*
X-0007163D01*
Y0016710D01*
X0034007Y-0031173D02*
X0033832D01*
X0033920Y-0030998D01*
X0033963D01*
Y-0031261D01*
X0033653Y-0031130D02*
X0033478D01*
X0033653Y-0031261D02*
Y-0030998D01*
X0033478Y-0031261D02*
Y-0030998D01*
X0033211Y-0031261D02*
Y-0030998D01*
X0033299D02*
X0033124D01*
X0032944Y-0031261D02*
Y-0030998D01*
X0032900Y-0031042D01*
X0032857Y-0031130D01*
X0032813Y-0031042D01*
X0032769Y-0030998D01*
Y-0031261D01*
X0035029Y-0032871D02*
X0035073Y-0032915D01*
X0035160D01*
X0035204Y-0032871D01*
Y-0032827D01*
X0035117Y-0032739D01*
X0035204Y-0032652D01*
X0035029D01*
X0034850Y-0032783D02*
X0034675D01*
X0034850Y-0032915D02*
Y-0032652D01*
X0034675Y-0032915D02*
Y-0032652D01*
X0034408Y-0032915D02*
Y-0032652D01*
X0034496D02*
X0034320D01*
X0034141Y-0032915D02*
Y-0032652D01*
X0034097Y-0032696D01*
X0034054Y-0032783D01*
X0034010Y-0032696D01*
X0033966Y-0032652D01*
Y-0032915D01*
X-0004119Y0016491D02*
X-0004076Y0016448D01*
X-0003988D01*
X-0003944Y0016491D01*
Y0016535D01*
X-0004032Y0016623D01*
X-0003944Y0016710D01*
X-0004119D01*
X-0004298Y0016448D02*
X-0004386D01*
X-0004342D02*
Y0016710D01*
X-0004386Y0016667D01*
X-0004762Y0016448D02*
Y0016710D01*
X-0004784Y0016448D02*
X-0004653D01*
X-0004609Y0016535D01*
Y0016623D01*
X-0004653Y0016710D01*
X-0004784D01*
X-0005007Y0016579D02*
X-0005138D01*
X-0004963Y0016448D02*
X-0005138D01*
Y0016710D01*
X-0004963D01*
X-0005317Y0016448D02*
X-0005470D01*
Y0016710D01*
X0031941Y-0032025D02*
X0031765D01*
X0031941Y-0031850D01*
Y-0031806D01*
X0031919Y-0031762D01*
X0031787D01*
X0031765Y-0031806D01*
X0031586Y-0031893D02*
X0031411D01*
X0031586Y-0032025D02*
Y-0031762D01*
X0031411Y-0032025D02*
Y-0031762D01*
X0031144Y-0032025D02*
Y-0031762D01*
X0031232D02*
X0031057D01*
X0030878Y-0032025D02*
Y-0031762D01*
X0030833Y-0031806D01*
X0030790Y-0031893D01*
X0030746Y-0031806D01*
X0030702Y-0031762D01*
Y-0032025D01*
X0033881Y-0031631D02*
X0033793D01*
X0033837D02*
Y-0031369D01*
X0033793Y-0031412D01*
X0033570Y-0031500D02*
X0033395D01*
X0033570Y-0031631D02*
Y-0031369D01*
X0033395Y-0031631D02*
Y-0031369D01*
X0033128Y-0031631D02*
Y-0031369D01*
X0033216D02*
X0033041D01*
X0032862Y-0031631D02*
Y-0031369D01*
X0032818Y-0031412D01*
X0032774Y-0031500D01*
X0032730Y-0031412D01*
X0032687Y-0031369D01*
Y-0031631D01*
X-0009128Y0015326D02*
X-0008996Y0015588D01*
X-0009171D01*
X-0009350D02*
Y0015369D01*
X-0009372Y0015326D01*
X-0009504D01*
X-0009526Y0015369D01*
Y0015588D01*
X0035084Y-0032056D02*
X0034997D01*
X0035041D02*
Y-0031794D01*
X0034997Y-0031837D01*
X0034774Y-0032056D02*
X0034687D01*
X0034730D02*
Y-0031794D01*
X0034687Y-0031837D01*
X0034464Y-0032056D02*
X0034376D01*
X0034420D02*
Y-0031794D01*
X0034376Y-0031837D01*
X0034154Y-0031794D02*
Y-0031881D01*
X0034066Y-0032056D01*
X0033978Y-0031881D01*
Y-0031794D01*
X0033624Y-0031925D02*
X0033755D01*
X0033799Y-0031881D01*
Y-0031837D01*
X0033755Y-0031794D01*
X0033624D01*
Y-0032056D01*
X0035920Y-0032758D02*
X0035877Y-0032802D01*
Y-0032889D01*
X0035920Y-0032933D01*
X0035965D01*
X0036052Y-0032845D01*
X0036139Y-0032933D01*
Y-0032758D01*
Y-0032579D02*
X0036052D01*
X0035877Y-0032491D01*
X0036052Y-0032404D01*
X0036139D01*
X0036008Y-0032049D02*
Y-0032180D01*
X0036052Y-0032224D01*
X0036096D01*
X0036139Y-0032180D01*
Y-0032049D01*
X0035877D01*
X-0016739Y0016448D02*
X-0016915D01*
X-0016739Y0016623D01*
Y0016667D01*
X-0016761Y0016710D01*
X-0016893D01*
X-0016915Y0016667D01*
X-0017094Y0016448D02*
X-0017181D01*
X-0017137D02*
Y0016710D01*
X-0017181Y0016667D01*
X-0017557Y0016448D02*
Y0016710D01*
X-0017579Y0016448D02*
X-0017448D01*
X-0017404Y0016535D01*
Y0016623D01*
X-0017448Y0016710D01*
X-0017579D01*
X-0017802Y0016579D02*
X-0017933D01*
X-0017758Y0016448D02*
X-0017933D01*
Y0016710D01*
X-0017758D01*
X-0018113Y0016448D02*
X-0018266D01*
Y0016710D01*
X0036270Y-0032408D02*
X0036533Y-0032539D01*
Y-0032364D01*
Y-0032185D02*
X0036446D01*
X0036270Y-0032097D01*
X0036446Y-0032010D01*
X0036533D01*
X0036402Y-0031656D02*
Y-0031787D01*
X0036446Y-0031831D01*
X0036489D01*
X0036533Y-0031787D01*
Y-0031656D01*
X0036270D01*
X0006826Y0016579D02*
X0006695D01*
X0006673Y0016623D01*
Y0016667D01*
X0006695Y0016710D01*
X0006826D01*
X0006848Y0016667D01*
Y0016623D01*
X0006760Y0016448D01*
X0006341D02*
Y0016710D01*
X0006319Y0016448D02*
X0006450D01*
X0006494Y0016535D01*
Y0016623D01*
X0006450Y0016710D01*
X0006319D01*
X0006095Y0016579D02*
X0005964D01*
X0006139Y0016448D02*
X0005964D01*
Y0016710D01*
X0006139D01*
X0005785Y0016448D02*
X0005632D01*
Y0016710D01*
X0035571Y-0032933D02*
Y-0032758D01*
X0035746Y-0032845D01*
Y-0032889D01*
X0035483D01*
X0035746Y-0032579D02*
X0035658D01*
X0035483Y-0032491D01*
X0035658Y-0032404D01*
X0035746D01*
X0035615Y-0032049D02*
Y-0032180D01*
X0035658Y-0032224D01*
X0035702D01*
X0035746Y-0032180D01*
Y-0032049D01*
X0035483D01*
X0035133Y-0032758D02*
X0035089Y-0032780D01*
Y-0032911D01*
X0035133Y-0032933D01*
X0035221D01*
X0035265Y-0032889D01*
Y-0032758D01*
X0035352D01*
Y-0032933D01*
Y-0032579D02*
X0035265D01*
X0035089Y-0032491D01*
X0035265Y-0032404D01*
X0035352D01*
X0035221Y-0032049D02*
Y-0032180D01*
X0035265Y-0032224D01*
X0035308D01*
X0035352Y-0032180D01*
Y-0032049D01*
X0035089D01*
X0001931Y0015369D02*
X0001953Y0015326D01*
X0002084D01*
X0002106Y0015369D01*
Y0015457D01*
X0002062Y0015501D01*
X0001931D01*
Y0015588D01*
X0002106D01*
X0001752D02*
Y0015369D01*
X0001730Y0015326D01*
X0001599D01*
X0001577Y0015369D01*
Y0015588D01*
X0033093Y-0032141D02*
X0033071Y-0032097D01*
X0032940D01*
X0032918Y-0032141D01*
Y-0032229D01*
X0032962Y-0032272D01*
X0033093D01*
Y-0032360D01*
X0032918D01*
X0033382Y-0032097D02*
X0033426Y-0032141D01*
X0033448Y-0032185D01*
Y-0032272D01*
X0033426Y-0032316D01*
X0033382Y-0032360D01*
X0033338D01*
X0033294Y-0032316D01*
X0033272Y-0032272D01*
Y-0032185D01*
X0033294Y-0032141D01*
X0033338Y-0032097D01*
X0033382D01*
X0033627D02*
X0033714D01*
X0033670D02*
Y-0032360D01*
X0033714Y-0032316D01*
X0033937Y-0032360D02*
Y-0032272D01*
X0034025Y-0032097D01*
X0034112Y-0032272D01*
Y-0032360D01*
X0034467Y-0032229D02*
X0034335D01*
X0034291Y-0032272D01*
Y-0032316D01*
X0034335Y-0032360D01*
X0034467D01*
Y-0032097D01*
X0036796Y-0032386D02*
Y-0032517D01*
X0036752Y-0032539D01*
X0036708D01*
X0036664Y-0032517D01*
Y-0032386D01*
X0036708Y-0032364D01*
X0036752D01*
X0036927Y-0032452D01*
Y-0032185D02*
X0036839D01*
X0036664Y-0032097D01*
X0036839Y-0032010D01*
X0036927D01*
X0036796Y-0031656D02*
Y-0031787D01*
X0036839Y-0031831D01*
X0036883D01*
X0036927Y-0031787D01*
Y-0031656D01*
X0036664D01*
X0016550Y0016579D02*
X0016572Y0016623D01*
Y0016667D01*
X0016550Y0016710D01*
X0016419D01*
X0016397Y0016667D01*
Y0016623D01*
X0016419Y0016579D01*
X0016550D01*
X0016572Y0016535D01*
Y0016491D01*
X0016550Y0016448D01*
X0016419D01*
X0016397Y0016491D01*
Y0016535D01*
X0016419Y0016579D01*
X0016065Y0016448D02*
Y0016710D01*
X0016043Y0016448D02*
X0016174D01*
X0016218Y0016535D01*
Y0016623D01*
X0016174Y0016710D01*
X0016043D01*
X0015820Y0016579D02*
X0015689D01*
X0015864Y0016448D02*
X0015689D01*
Y0016710D01*
X0015864D01*
X0015509Y0016448D02*
X0015356D01*
Y0016710D01*
X0017819Y0016448D02*
X0017950Y0016710D01*
X0017775D01*
X0017443Y0016448D02*
Y0016710D01*
X0017421Y0016448D02*
X0017552D01*
X0017596Y0016535D01*
Y0016623D01*
X0017552Y0016710D01*
X0017421D01*
X0017198Y0016579D02*
X0017067D01*
X0017242Y0016448D02*
X0017067D01*
Y0016710D01*
X0017242D01*
X0016887Y0016448D02*
X0016734D01*
Y0016710D01*
X0013189Y0015413D02*
X0013014D01*
X0013101Y0015588D01*
X0013145D01*
Y0015326D01*
X0012835Y0015588D02*
Y0015369D01*
X0012813Y0015326D01*
X0012681D01*
X0012659Y0015369D01*
Y0015588D01*
X0062198Y0034219D02*
X0062154Y0034306D01*
X0061892D01*
X0061848Y0034219D01*
Y0034131D01*
X0061892Y0034044D01*
X0062154D01*
X0062198Y0033957D01*
Y0033869D01*
X0062154Y0033781D01*
X0061892D01*
X0061848Y0033869D01*
X0061341Y0033781D02*
X0061297Y0033869D01*
Y0034219D01*
X0061341Y0034306D01*
X0061603D01*
X0061647Y0034219D01*
Y0033869D01*
X0061603Y0033781D01*
X0061341D01*
X0061096D02*
Y0034306D01*
X0061008Y0034219D01*
X0060921Y0034044D01*
X0060833Y0034219D01*
X0060746Y0034306D01*
Y0033781D01*
X0060545D02*
X0060283Y0034306D01*
X0060545D02*
X0060283Y0033781D01*
X0059290D02*
Y0034306D01*
X0059202Y0034219D01*
X0059115Y0034044D01*
X0059027Y0034219D01*
X0058940Y0034306D01*
Y0033781D01*
X0058432D02*
X0058389Y0033869D01*
Y0034219D01*
X0058432Y0034306D01*
X0058694D01*
X0058739Y0034219D01*
Y0033869D01*
X0058694Y0033781D01*
X0058432D01*
X0058056Y0034044D02*
X0058187Y0033781D01*
X0057837Y0034044D02*
X0058100D01*
X0058187Y0034131D01*
Y0034219D01*
X0058100Y0034306D01*
X0057837D01*
Y0033781D01*
X0057548Y0034044D02*
X0057286D01*
Y0033781D02*
Y0034306D01*
X0057636D01*
X0056337D02*
Y0033781D01*
X0056249Y0033869D01*
X0056074Y0034219D01*
X0055987Y0034306D01*
Y0033781D01*
X0055480D02*
X0055436Y0033869D01*
Y0034219D01*
X0055480Y0034306D01*
X0055742D01*
X0055786Y0034219D01*
Y0033869D01*
X0055742Y0033781D01*
X0055480D01*
X0055235D02*
X0055060D01*
X0055147D02*
Y0034306D01*
X0055235D02*
X0055060D01*
X0054596Y0033781D02*
Y0034306D01*
X0054771D02*
X0054421D01*
X0054220Y0033869D02*
X0054176Y0033781D01*
X0053914D01*
X0053870Y0033869D01*
Y0034219D01*
X0053914Y0034306D01*
X0054176D01*
X0054220Y0034219D01*
X0053669Y0034306D02*
Y0033869D01*
X0053625Y0033781D01*
X0053363D01*
X0053319Y0033869D01*
Y0034306D01*
X0052986Y0034044D02*
X0053118Y0033781D01*
X0052768Y0034044D02*
X0053030D01*
X0053118Y0034131D01*
Y0034219D01*
X0053030Y0034306D01*
X0052768D01*
Y0033781D01*
X0052391D02*
Y0034306D01*
X0052567D02*
X0052217D01*
X0052015Y0034219D02*
X0051971Y0034306D01*
X0051709D01*
X0051665Y0034219D01*
Y0034131D01*
X0051709Y0034044D01*
X0051971D01*
X0052015Y0033957D01*
Y0033869D01*
X0051971Y0033781D01*
X0051709D01*
X0051665Y0033869D01*
X0051464Y0034306D02*
Y0033781D01*
X0051376Y0033869D01*
X0051202Y0034219D01*
X0051114Y0034306D01*
Y0033781D01*
X0050913D02*
X0050738D01*
X0050826D02*
Y0034306D01*
X0050913D02*
X0050738D01*
X0049702Y0034044D02*
X0049352D01*
X0048096Y0033781D02*
Y0034306D01*
X0048052Y0033781D02*
X0048315D01*
X0048402Y0033957D01*
Y0034131D01*
X0048315Y0034306D01*
X0048052D01*
X0047763Y0034044D02*
X0047501D01*
X0047851Y0033781D02*
X0047501D01*
Y0034306D01*
X0047851D01*
X0047300Y0034044D02*
X0046950D01*
X0047300Y0033781D02*
Y0034306D01*
X0046950Y0033781D02*
Y0034306D01*
X0046574Y0033781D02*
Y0034306D01*
X0046749D02*
X0046399D01*
X0046022Y0034044D02*
X0046198D01*
Y0033869D01*
X0046154Y0033781D01*
X0045891D01*
X0045848Y0033869D01*
Y0034219D01*
X0045891Y0034306D01*
X0046154D01*
X0046198Y0034219D01*
X0045646Y0034306D02*
Y0033781D01*
X0045559Y0033869D01*
X0045384Y0034219D01*
X0045296Y0034306D01*
Y0033781D01*
X0045007Y0034044D02*
X0044745D01*
X0045095Y0033781D02*
X0044745D01*
Y0034306D01*
X0045095D01*
X0044544Y0033781D02*
X0044238D01*
Y0034306D01*
X0043289Y0034044D02*
X0042939D01*
X0043289Y0033781D02*
Y0034306D01*
X0042939Y0033781D02*
Y0034306D01*
X0042738Y0033869D02*
X0042694Y0033781D01*
X0042431D01*
X0042388Y0033869D01*
Y0034219D01*
X0042431Y0034306D01*
X0042694D01*
X0042738Y0034219D01*
X0042011Y0033781D02*
Y0034306D01*
X0042187D02*
X0041837D01*
X0041635Y0033957D02*
X0041285D01*
X0041635Y0033781D02*
Y0034044D01*
X0041504Y0034306D01*
X0041417D01*
X0041285Y0034044D01*
Y0033781D01*
X0041084D02*
Y0034306D01*
X0040996Y0034219D01*
X0040909Y0034044D01*
X0040822Y0034219D01*
X0040734Y0034306D01*
Y0033781D01*
X0039697Y0034044D02*
X0039435D01*
X0039785Y0033781D02*
X0039435D01*
Y0034306D01*
X0039785D01*
X0038928Y0033781D02*
Y0034306D01*
X0038884Y0033781D02*
X0039146D01*
X0039234Y0033869D01*
Y0033957D01*
X0039190Y0034044D01*
X0038928D02*
X0039190D01*
X0039234Y0034131D01*
Y0034219D01*
X0039146Y0034306D01*
X0038884D01*
X0037628Y0033781D02*
X0037585Y0033869D01*
Y0034219D01*
X0037628Y0034306D01*
X0037891D01*
X0037935Y0034219D01*
Y0033869D01*
X0037891Y0033781D01*
X0037628D01*
X0037208D02*
Y0034306D01*
X0037383D02*
X0037033D01*
X0035778Y0033781D02*
Y0034306D01*
X0035734Y0033781D02*
X0035996D01*
X0036084Y0033957D01*
Y0034131D01*
X0035996Y0034306D01*
X0035734D01*
X0035445Y0034044D02*
X0035183D01*
X0035533Y0033781D02*
X0035183D01*
Y0034306D01*
X0035533D01*
X0034894Y0034044D02*
X0034632D01*
X0034982Y0033781D02*
X0034632D01*
Y0034306D01*
X0034982D01*
X0034431D02*
Y0033781D01*
X0034343Y0033869D01*
X0034168Y0034219D01*
X0034081Y0034306D01*
Y0033781D01*
X0032956D02*
Y0034306D01*
X0033131D02*
X0032781D01*
X0032537Y0034219D02*
X0032580Y0034306D01*
X0032161D02*
Y0033781D01*
X0032073Y0033869D01*
X0031898Y0034219D01*
X0031811Y0034306D01*
Y0033781D01*
X0031303D02*
X0031259Y0033869D01*
Y0034219D01*
X0031303Y0034306D01*
X0031565D01*
X0031609Y0034219D01*
Y0033869D01*
X0031565Y0033781D01*
X0031303D01*
X0030752D02*
Y0034306D01*
X0030708Y0033781D02*
X0030970D01*
X0031058Y0033957D01*
Y0034131D01*
X0030970Y0034306D01*
X0030708D01*
X0029759Y0034219D02*
X0029715Y0034306D01*
X0029453D01*
X0029409Y0034219D01*
Y0034131D01*
X0029453Y0034044D01*
X0029715D01*
X0029759Y0033957D01*
Y0033869D01*
X0029715Y0033781D01*
X0029453D01*
X0029409Y0033869D01*
X0029208Y0033781D02*
X0028945Y0034044D01*
X0029208Y0034306D01*
X0028858D02*
Y0033781D01*
X0028657Y0033869D02*
X0028613Y0033781D01*
X0028350D01*
X0028307Y0033869D01*
Y0034219D01*
X0028350Y0034306D01*
X0028613D01*
X0028657Y0034219D01*
X0027799Y0033781D02*
X0027756Y0033869D01*
Y0034219D01*
X0027799Y0034306D01*
X0028061D01*
X0028106Y0034219D01*
Y0033869D01*
X0028061Y0033781D01*
X0027799D01*
X0027554D02*
X0027248D01*
Y0034306D01*
X0027047Y0033869D02*
X0027003Y0033781D01*
X0026741D01*
X0026697Y0033869D01*
Y0034219D01*
X0026741Y0034306D01*
X0027003D01*
X0027047Y0034219D01*
X0035019Y-0031781D02*
X0034975Y-0031737D01*
X0034953Y-0031693D01*
Y-0031606D01*
X0034975Y-0031562D01*
X0035019Y-0031518D01*
X0035063D01*
X0035106Y-0031562D01*
X0035128Y-0031606D01*
Y-0031693D01*
X0035106Y-0031737D01*
X0035063Y-0031781D01*
X0035019D01*
X0034774D02*
X0034687D01*
X0034730D02*
Y-0031518D01*
X0034687Y-0031562D01*
X0034464Y-0031781D02*
X0034376D01*
X0034420D02*
Y-0031518D01*
X0034376Y-0031562D01*
X0034154Y-0031518D02*
Y-0031606D01*
X0034066Y-0031781D01*
X0033978Y-0031606D01*
Y-0031518D01*
X0033624Y-0031649D02*
X0033755D01*
X0033799Y-0031606D01*
Y-0031562D01*
X0033755Y-0031518D01*
X0033624D01*
Y-0031781D01*
X0035615Y-0032517D02*
Y-0032386D01*
X0035658Y-0032364D01*
X0035702D01*
X0035746Y-0032386D01*
Y-0032517D01*
X0035702Y-0032539D01*
X0035658D01*
X0035483Y-0032452D01*
X0035746Y-0032185D02*
X0035658D01*
X0035483Y-0032097D01*
X0035658Y-0032010D01*
X0035746D01*
X0035615Y-0031656D02*
Y-0031787D01*
X0035658Y-0031831D01*
X0035702D01*
X0035746Y-0031787D01*
Y-0031656D01*
X0035483D01*
X0005356Y0016448D02*
X0005312Y0016491D01*
X0005290Y0016535D01*
Y0016623D01*
X0005312Y0016667D01*
X0005356Y0016710D01*
X0005400D01*
X0005443Y0016667D01*
X0005465Y0016623D01*
Y0016535D01*
X0005443Y0016491D01*
X0005400Y0016448D01*
X0005356D01*
X0005111D02*
X0005024D01*
X0005067D02*
Y0016710D01*
X0005024Y0016667D01*
X0004648Y0016448D02*
Y0016710D01*
X0004626Y0016448D02*
X0004757D01*
X0004801Y0016535D01*
Y0016623D01*
X0004757Y0016710D01*
X0004626D01*
X0004402Y0016579D02*
X0004271D01*
X0004446Y0016448D02*
X0004271D01*
Y0016710D01*
X0004446D01*
X0004092Y0016448D02*
X0003939D01*
Y0016710D01*
X-0015134Y0005345D02*
X-0015002Y0005608D01*
X-0015178D01*
X-0015357Y0005345D02*
X-0015532D01*
X-0015357Y0005520D01*
Y0005564D01*
X-0015379Y0005608D01*
X-0015510D01*
X-0015532Y0005564D01*
X-0015864Y0005345D02*
Y0005608D01*
X-0015886Y0005345D02*
X-0015755D01*
X-0015711Y0005433D01*
Y0005520D01*
X-0015755Y0005608D01*
X-0015886D01*
X-0016109Y0005477D02*
X-0016241D01*
X-0016065Y0005345D02*
X-0016241D01*
Y0005608D01*
X-0016065D01*
X-0016420Y0005345D02*
X-0016573D01*
Y0005608D01*
X-0004430Y0027594D02*
X-0004407Y0027550D01*
X-0004276D01*
X-0004254Y0027594D01*
Y0027681D01*
X-0004298Y0027725D01*
X-0004430D01*
Y0027813D01*
X-0004254D01*
X-0004762Y0027550D02*
Y0027813D01*
X-0004784Y0027550D02*
X-0004653D01*
X-0004609Y0027638D01*
Y0027725D01*
X-0004653Y0027813D01*
X-0004784D01*
X-0005007Y0027681D02*
X-0005138D01*
X-0004963Y0027550D02*
X-0005138D01*
Y0027813D01*
X-0004963D01*
X-0005317Y0027550D02*
X-0005470D01*
Y0027813D01*
X0035546Y-0033001D02*
X0035371D01*
X0035546Y-0032826D01*
Y-0032782D01*
X0035524Y-0032739D01*
X0035393D01*
X0035371Y-0032782D01*
X0035017Y-0032957D02*
X0035039Y-0033001D01*
X0035170D01*
X0035192Y-0032957D01*
Y-0032870D01*
X0035148Y-0032826D01*
X0035017D01*
Y-0032739D01*
X0035192D01*
X0034838Y-0033001D02*
X0034750D01*
X0034794D02*
Y-0032739D01*
X0034750Y-0032782D01*
X0034528Y-0032739D02*
Y-0032826D01*
X0034440Y-0033001D01*
X0034352Y-0032826D01*
Y-0032739D01*
X0033998Y-0032870D02*
X0034129D01*
X0034173Y-0032826D01*
Y-0032782D01*
X0034129Y-0032739D01*
X0033998D01*
Y-0033001D01*
X-0009171Y0026491D02*
X-0009128Y0026448D01*
X-0009040D01*
X-0008996Y0026491D01*
Y0026535D01*
X-0009084Y0026623D01*
X-0008996Y0026710D01*
X-0009171D01*
X-0009350D02*
Y0026491D01*
X-0009372Y0026448D01*
X-0009504D01*
X-0009526Y0026491D01*
Y0026710D01*
X0034057Y-0033513D02*
X0034188Y-0033250D01*
X0034013D01*
X0033724Y-0033513D02*
X0033681Y-0033469D01*
X0033659Y-0033425D01*
Y-0033338D01*
X0033681Y-0033294D01*
X0033724Y-0033250D01*
X0033768D01*
X0033812Y-0033294D01*
X0033834Y-0033338D01*
Y-0033425D01*
X0033812Y-0033469D01*
X0033768Y-0033513D01*
X0033724D01*
X0033480D02*
X0033392D01*
X0033436D02*
Y-0033250D01*
X0033392Y-0033294D01*
X0033169Y-0033250D02*
Y-0033338D01*
X0033081Y-0033513D01*
X0032994Y-0033338D01*
Y-0033250D01*
X0032640Y-0033381D02*
X0032771D01*
X0032815Y-0033338D01*
Y-0033294D01*
X0032771Y-0033250D01*
X0032640D01*
Y-0033513D01*
X-0005785Y0027681D02*
X-0005654D01*
X-0005632Y0027638D01*
Y0027594D01*
X-0005654Y0027550D01*
X-0005785D01*
X-0005807Y0027594D01*
Y0027638D01*
X-0005720Y0027813D01*
X-0006140Y0027550D02*
Y0027813D01*
X-0006162Y0027550D02*
X-0006031D01*
X-0005987Y0027638D01*
Y0027725D01*
X-0006031Y0027813D01*
X-0006162D01*
X-0006385Y0027681D02*
X-0006516D01*
X-0006341Y0027550D02*
X-0006516D01*
Y0027813D01*
X-0006341D01*
X-0006695Y0027550D02*
X-0006848D01*
Y0027813D01*
X0064479Y0021999D02*
Y0022261D01*
X0064567D02*
X0064392D01*
X0064213Y0021999D02*
Y0022261D01*
X0064169Y0022218D01*
X0064125Y0022130D01*
X0064081Y0022218D01*
X0064037Y0022261D01*
Y0021999D01*
X0063858Y0022218D02*
X0063836Y0022261D01*
X0063705D01*
X0063683Y0022218D01*
Y0022174D01*
X0063705Y0022130D01*
X0063836D01*
X0063858Y0022087D01*
Y0022043D01*
X0063836Y0021999D01*
X0063705D01*
X0063683Y0022043D01*
X-0015532Y0027574D02*
X-0015488Y0027530D01*
X-0015401D01*
X-0015357Y0027574D01*
Y0027618D01*
X-0015444Y0027706D01*
X-0015357Y0027793D01*
X-0015532D01*
X-0015864Y0027530D02*
Y0027793D01*
X-0015886Y0027530D02*
X-0015755D01*
X-0015711Y0027618D01*
Y0027706D01*
X-0015755Y0027793D01*
X-0015886D01*
X-0016109Y0027662D02*
X-0016241D01*
X-0016065Y0027530D02*
X-0016241D01*
Y0027793D01*
X-0016065D01*
X-0016420Y0027530D02*
X-0016573D01*
Y0027793D01*
X0074228Y0022918D02*
X0074359D01*
X0074404Y0022961D01*
Y0023005D01*
X0074359Y0023049D01*
X0074228D01*
Y0022786D01*
X0073896D02*
X0073874Y0022830D01*
Y0023005D01*
X0073896Y0023049D01*
X0074027D01*
X0074049Y0023005D01*
Y0022830D01*
X0074027Y0022786D01*
X0073896D01*
X0073607D02*
Y0023049D01*
X0073695D02*
X0073520D01*
X0072844Y0022786D02*
X0072888Y0022874D01*
Y0022961D01*
X0072844Y0023049D01*
X0072533Y0022786D02*
Y0023049D01*
X0072621D02*
X0072446D01*
X0072267D02*
Y0022786D01*
X0072223Y0022830D01*
X0072135Y0023005D01*
X0072092Y0023049D01*
Y0022786D01*
X0071869Y0022918D02*
X0071737D01*
X0071913Y0022786D02*
X0071737D01*
Y0023049D01*
X0071913D01*
X0071405Y0022786D02*
Y0023049D01*
X0071383Y0022786D02*
X0071514D01*
X0071558Y0022874D01*
Y0022961D01*
X0071514Y0023049D01*
X0071383D01*
X0071204Y0022786D02*
X0071117D01*
X0071160D02*
Y0023049D01*
X0071204D02*
X0071117D01*
X0070894Y0022786D02*
X0070850Y0022874D01*
Y0022961D01*
X0070894Y0023049D01*
X0070131D02*
Y0022786D01*
X0070087Y0022830D01*
X0069999Y0023005D01*
X0069956Y0023049D01*
Y0022786D01*
X0069732Y0022918D02*
X0069601D01*
X0069776Y0022786D02*
X0069601D01*
Y0023049D01*
X0069776D01*
X0069378Y0022918D02*
X0069247D01*
X0069422Y0022786D02*
X0069247D01*
Y0023049D01*
X0069422D01*
X0069002Y0022918D02*
X0069068Y0022786D01*
X0068893Y0022918D02*
X0069024D01*
X0069068Y0022961D01*
Y0023005D01*
X0069024Y0023049D01*
X0068893D01*
Y0022786D01*
X0068713Y0022830D02*
X0068691Y0022786D01*
X0068560D01*
X0068538Y0022830D01*
Y0023005D01*
X0068560Y0023049D01*
X0068691D01*
X0068713Y0023005D01*
X0068359D02*
X0068337Y0023049D01*
X0068206D01*
X0068184Y0023005D01*
Y0022961D01*
X0068206Y0022918D01*
X0068337D01*
X0068359Y0022874D01*
Y0022830D01*
X0068337Y0022786D01*
X0068206D01*
X0068184Y0022830D01*
X0068005Y0022786D02*
X0067873Y0022918D01*
X0068005Y0023049D01*
X0067830D02*
Y0022786D01*
X0067650D02*
X0067497D01*
Y0023049D01*
X0067318Y0022786D02*
X0067231D01*
X0067274D02*
Y0023049D01*
X0067318D02*
X0067231D01*
X0067008Y0023005D02*
X0066986Y0023049D01*
X0066855D01*
X0066833Y0023005D01*
Y0022961D01*
X0066855Y0022918D01*
X0066986D01*
X0067008Y0022874D01*
Y0022830D01*
X0066986Y0022786D01*
X0066855D01*
X0066833Y0022830D01*
X-0020098Y0026428D02*
X-0020274D01*
X-0020098Y0026603D01*
Y0026647D01*
X-0020120Y0026691D01*
X-0020252D01*
X-0020274Y0026647D01*
X-0020453Y0026691D02*
Y0026472D01*
X-0020475Y0026428D01*
X-0020606D01*
X-0020628Y0026472D01*
Y0026691D01*
X0033312Y-0031782D02*
X0033487D01*
X0033312Y-0031957D01*
Y-0032001D01*
X0033334Y-0032045D01*
X0033465D01*
X0033487Y-0032001D01*
X0033776Y-0031782D02*
X0033819Y-0031826D01*
X0033841Y-0031870D01*
Y-0031957D01*
X0033819Y-0032001D01*
X0033776Y-0032045D01*
X0033732D01*
X0033688Y-0032001D01*
X0033666Y-0031957D01*
Y-0031870D01*
X0033688Y-0031826D01*
X0033732Y-0031782D01*
X0033776D01*
X0034020D02*
X0034108D01*
X0034064D02*
Y-0032045D01*
X0034108Y-0032001D01*
X0034331Y-0032045D02*
Y-0031957D01*
X0034419Y-0031782D01*
X0034506Y-0031957D01*
Y-0032045D01*
X0034860Y-0031914D02*
X0034729D01*
X0034685Y-0031957D01*
Y-0032001D01*
X0034729Y-0032045D01*
X0034860D01*
Y-0031782D01*
X-0016735Y0027618D02*
X-0016910D01*
X-0016822Y0027793D01*
X-0016779D01*
Y0027530D01*
X-0017242D02*
Y0027793D01*
X-0017264Y0027530D02*
X-0017133D01*
X-0017089Y0027618D01*
Y0027706D01*
X-0017133Y0027793D01*
X-0017264D01*
X-0017487Y0027662D02*
X-0017619D01*
X-0017443Y0027530D02*
X-0017619D01*
Y0027793D01*
X-0017443D01*
X-0017798Y0027530D02*
X-0017951D01*
Y0027793D01*
X0002062Y0026448D02*
X0001975D01*
X0002019D02*
Y0026710D01*
X0001975Y0026667D01*
X0001752Y0026710D02*
Y0026491D01*
X0001730Y0026448D01*
X0001599D01*
X0001577Y0026491D01*
Y0026710D01*
X0018130Y0027594D02*
X0018173Y0027550D01*
X0018261D01*
X0018305Y0027594D01*
Y0027638D01*
X0018217Y0027725D01*
X0018305Y0027813D01*
X0018130D01*
X0017775Y0027594D02*
X0017819Y0027550D01*
X0017906D01*
X0017950Y0027594D01*
Y0027638D01*
X0017863Y0027725D01*
X0017950Y0027813D01*
X0017775D01*
X0017443Y0027550D02*
Y0027813D01*
X0017421Y0027550D02*
X0017552D01*
X0017596Y0027638D01*
Y0027725D01*
X0017552Y0027813D01*
X0017421D01*
X0017198Y0027681D02*
X0017067D01*
X0017242Y0027550D02*
X0017067D01*
Y0027813D01*
X0017242D01*
X0016887Y0027550D02*
X0016734D01*
Y0027813D01*
X0075080Y0022130D02*
X0075211D01*
X0075255Y0022174D01*
Y0022218D01*
X0075211Y0022261D01*
X0075080D01*
Y0021999D01*
X0074747D02*
X0074725Y0022043D01*
Y0022218D01*
X0074747Y0022261D01*
X0074878D01*
X0074900Y0022218D01*
Y0022043D01*
X0074878Y0021999D01*
X0074747D01*
X0074458D02*
Y0022261D01*
X0074546D02*
X0074371D01*
X0073695Y0021999D02*
X0073739Y0022087D01*
Y0022174D01*
X0073695Y0022261D01*
X0073385Y0021999D02*
Y0022261D01*
X0073472D02*
X0073297D01*
X0073118Y0022218D02*
X0073096Y0022261D01*
X0072965D01*
X0072943Y0022218D01*
Y0022174D01*
X0072965Y0022130D01*
X0073096D01*
X0073118Y0022087D01*
Y0022043D01*
X0073096Y0021999D01*
X0072965D01*
X0072943Y0022043D01*
X0072764Y0021999D02*
X0072676D01*
X0072720D02*
Y0022261D01*
X0072764D02*
X0072676D01*
X0072454Y0022218D02*
X0072431Y0022261D01*
X0072300D01*
X0072278Y0022218D01*
Y0022174D01*
X0072300Y0022130D01*
X0072431D01*
X0072454Y0022087D01*
Y0022043D01*
X0072431Y0021999D01*
X0072300D01*
X0072278Y0022043D01*
X0072055Y0022130D02*
X0071924D01*
X0072099Y0021999D02*
X0071924D01*
Y0022261D01*
X0072099D01*
X0071679Y0022130D02*
X0071745Y0021999D01*
X0071570Y0022130D02*
X0071701D01*
X0071745Y0022174D01*
Y0022218D01*
X0071701Y0022261D01*
X0071570D01*
Y0021999D01*
X0071391D02*
X0071347Y0022087D01*
Y0022174D01*
X0071391Y0022261D01*
X0070628Y0021999D02*
X0070496Y0022130D01*
X0070628Y0022261D01*
X0070452D02*
Y0021999D01*
X0070273Y0022218D02*
X0070251Y0022261D01*
X0070120D01*
X0070098Y0022218D01*
Y0022174D01*
X0070120Y0022130D01*
X0070251D01*
X0070273Y0022087D01*
Y0022043D01*
X0070251Y0021999D01*
X0070120D01*
X0070098Y0022043D01*
X0069919Y0022087D02*
X0069744D01*
X0069919Y0021999D02*
Y0022130D01*
X0069853Y0022261D01*
X0069809D01*
X0069744Y0022130D01*
Y0021999D01*
X0069565D02*
Y0022261D01*
X0069520Y0022218D01*
X0069477Y0022130D01*
X0069433Y0022218D01*
X0069389Y0022261D01*
Y0021999D01*
X0068692Y0022130D02*
X0068757Y0021999D01*
X0068582Y0022130D02*
X0068713D01*
X0068757Y0022174D01*
Y0022218D01*
X0068713Y0022261D01*
X0068582D01*
Y0021999D01*
X0068359Y0022130D02*
X0068228D01*
X0068403Y0021999D02*
X0068228D01*
Y0022261D01*
X0068403D01*
X0067896Y0021999D02*
Y0022261D01*
X0067874Y0021999D02*
X0068005D01*
X0068049Y0022087D01*
Y0022174D01*
X0068005Y0022261D01*
X0067874D01*
X0067694Y0021999D02*
X0067541D01*
Y0022261D01*
X0067209Y0021999D02*
X0067187Y0022043D01*
Y0022218D01*
X0067209Y0022261D01*
X0067340D01*
X0067362Y0022218D01*
Y0022043D01*
X0067340Y0021999D01*
X0067209D01*
X0067008Y0022218D02*
X0066986Y0022261D01*
X0066855D01*
X0066833Y0022218D01*
Y0022174D01*
X0066855Y0022130D01*
X0066986D01*
X0067008Y0022087D01*
Y0022043D01*
X0066986Y0021999D01*
X0066855D01*
X0066833Y0022043D01*
X0006804Y0027550D02*
X0006717D01*
X0006760D02*
Y0027813D01*
X0006717Y0027769D01*
X0006341Y0027550D02*
Y0027813D01*
X0006319Y0027550D02*
X0006450D01*
X0006494Y0027638D01*
Y0027725D01*
X0006450Y0027813D01*
X0006319D01*
X0006095Y0027681D02*
X0005964D01*
X0006139Y0027550D02*
X0005964D01*
Y0027813D01*
X0006139D01*
X0005785Y0027550D02*
X0005632D01*
Y0027813D01*
X0005450Y0027550D02*
X0005275D01*
X0005450Y0027725D01*
Y0027769D01*
X0005428Y0027813D01*
X0005297D01*
X0005275Y0027769D01*
X0004943Y0027550D02*
Y0027813D01*
X0004921Y0027550D02*
X0005052D01*
X0005096Y0027638D01*
Y0027725D01*
X0005052Y0027813D01*
X0004921D01*
X0004698Y0027681D02*
X0004567D01*
X0004742Y0027550D02*
X0004567D01*
Y0027813D01*
X0004742D01*
X0004387Y0027550D02*
X0004234D01*
Y0027813D01*
X-0009575Y-0035228D02*
X-0007563D01*
Y-0034205D01*
X-0009575D01*
Y-0035228D01*
X0017343Y0026791D02*
Y0027303D01*
X0015965D02*
Y0026791D01*
X0012677Y0026280D02*
X0020630D01*
Y0018327D01*
X0012677D01*
Y0026280D01*
X0012913D02*
X0012677Y0026043D01*
X-0017343Y0005098D02*
Y0004587D01*
X-0015965D02*
Y0005098D01*
X-0020630Y0004075D02*
X-0012677D01*
Y-0003878D01*
X-0020630D01*
Y0004075D01*
X-0020394D02*
X-0020630Y0003839D01*
X-0006240Y0005098D02*
Y0004587D01*
X-0004862D02*
Y0005098D01*
X-0009528Y0004075D02*
X-0001575D01*
Y-0003878D01*
X-0009528D01*
Y0004075D01*
X-0009291D02*
X-0009528Y0003839D01*
X0004862Y0005098D02*
Y0004587D01*
X0006240D02*
Y0005098D01*
X0001575Y0004075D02*
X0009528D01*
Y-0003878D01*
X0001575D01*
Y0004075D01*
X0001811D02*
X0001575Y0003839D01*
X0015965Y0005098D02*
Y0004587D01*
X0017343D02*
Y0005098D01*
X0012677Y0004075D02*
X0020630D01*
Y-0003878D01*
X0012677D01*
Y0004075D01*
X0012913D02*
X0012677Y0003839D01*
X0004862Y-0006004D02*
Y-0006516D01*
X0006240D02*
Y-0006004D01*
X0001575Y-0007028D02*
X0009528D01*
Y-0014980D01*
X0001575D01*
Y-0007028D01*
X0001811D02*
X0001575Y-0007264D01*
X-0017343Y-0006004D02*
Y-0006516D01*
X-0023622Y0029134D02*
X-0022343D01*
X-0019390Y0032087D01*
X-0017815D01*
Y0031496D01*
X-0008031D01*
Y0035433D01*
X0008031D01*
Y0031457D01*
X0017953D01*
Y0032047D01*
X0019528D01*
X0022441Y0029134D01*
X0023622D01*
Y-0029134D01*
X0022244D01*
X0017244Y-0034134D01*
Y-0035433D01*
X-0017323D01*
Y-0034252D01*
X-0022441Y-0029134D01*
X-0023622D01*
Y0029134D01*
X-0015965Y-0006516D02*
Y-0006004D01*
X0023622Y0035039D02*
Y0035827D01*
X0023228Y0035433D02*
X0024016D01*
X0023622Y0035039D02*
Y0035827D01*
X0023228Y0035433D02*
X0024016D01*
X-0020630Y-0007028D02*
X-0012677D01*
Y-0014980D01*
X-0020630D01*
Y-0007028D01*
X-0020394D02*
X-0020630Y-0007264D01*
X-0006240Y-0006004D02*
Y-0006516D01*
X-0004862D02*
Y-0006004D01*
X-0009528Y-0007028D02*
X-0001575D01*
Y-0014980D01*
X-0009528D01*
Y-0007028D01*
X-0009291D02*
X-0009528Y-0007264D01*
X0015965Y-0006004D02*
Y-0006516D01*
X0017343D02*
Y-0006004D01*
X0012677Y-0007028D02*
X0020630D01*
Y-0014980D01*
X0012677D01*
Y-0007028D01*
X0012913D02*
X0012677Y-0007264D01*
X-0017343Y0016201D02*
Y0015689D01*
X-0015965D02*
Y0016201D01*
X-0020630Y0015177D02*
X-0012677D01*
Y0007224D01*
X-0020630D01*
Y0015177D01*
X-0020394D02*
X-0020630Y0014941D01*
X-0006240Y0016201D02*
Y0015689D01*
X-0004862D02*
Y0016201D01*
X-0009528Y0015177D02*
X-0001575D01*
Y0007224D01*
X-0009528D01*
Y0015177D01*
X-0009291D02*
X-0009528Y0014941D01*
X0004862Y0016201D02*
Y0015689D01*
X0006240D02*
Y0016201D01*
X0001575Y0015177D02*
X0009528D01*
Y0007224D01*
X0001575D01*
Y0015177D01*
X0001811D02*
X0001575Y0014941D01*
X0015965Y0016201D02*
Y0015689D01*
X0017343D02*
Y0016201D01*
X0012677Y0015177D02*
X0020630D01*
Y0007224D01*
X0012677D01*
Y0015177D01*
X0012913D02*
X0012677Y0014941D01*
X-0006240Y0027303D02*
Y0026791D01*
X-0004862D02*
Y0027303D01*
X-0009528Y0026280D02*
X-0001575D01*
Y0018327D01*
X-0009528D01*
Y0026280D01*
X-0009291D02*
X-0009528Y0026043D01*
X-0017343Y0027303D02*
Y0026791D01*
X-0015965D02*
Y0027303D01*
X-0020630Y0026280D02*
X-0012677D01*
Y0018327D01*
X-0020630D01*
Y0026280D01*
X-0020394D02*
X-0020630Y0026043D01*
X0001575Y0026280D02*
X0009528D01*
Y0018327D01*
X0001575D01*
Y0026280D01*
X0001811D02*
X0001575Y0026043D01*
X-0023622Y0029134D02*
X-0022343D01*
X-0019390Y0032087D01*
X-0017815D01*
Y0031496D01*
X-0008031D01*
Y0035433D01*
X0008031D01*
Y0031457D01*
X0017953D01*
Y0032047D01*
X0019528D01*
X0022441Y0029134D01*
X0023622D01*
Y-0029134D01*
X0022244D01*
X0017244Y-0034134D01*
Y-0035433D01*
X-0017323D01*
Y-0034252D01*
X-0022441Y-0029134D01*
X-0023622D01*
Y0029134D01*
Y-0035807D02*
Y-0035020D01*
X-0024016Y-0035413D02*
X-0023228D01*
X-0023622Y-0035807D02*
Y-0035020D01*
X-0024016Y-0035413D02*
X-0023228D01*
X0023622Y-0035807D02*
Y-0035020D01*
X0023228Y-0035413D02*
X0024016D01*
X0023622Y-0035807D02*
Y-0035020D01*
X0023228Y-0035413D02*
X0024016D01*
X0006240Y0026791D02*
Y0027303D01*
X0004862D02*
Y0026791D01*
G01X0012283Y0026555D02*
G03X0012401Y0026673I0000000J0000118D01*
G01X0012165D02*
G03X0012283Y0026555I0000118J0000000D01*
Y0026792D02*
G03X0012164Y0026673I0000000J0000119D01*
G01X0012402D02*
G03X0012283Y0026792I0000119J0000000D01*
G01X-0021024Y0004351D02*
G03X-0020906Y0004469I0000000J0000118D01*
G01X-0021142D02*
G03X-0021024Y0004351I0000118J0000000D01*
Y0004587D02*
G03X-0021142Y0004469I0000000J0000118D01*
G01X-0020906D02*
G03X-0021024Y0004587I0000118J0000000D01*
G01X-0009921Y0004351D02*
G03X-0009803Y0004469I0000000J0000118D01*
G01X-0010039D02*
G03X-0009921Y0004351I0000118J0000000D01*
Y0004587D02*
G03X-0010039Y0004469I0000000J0000118D01*
G01X-0009803D02*
G03X-0009921Y0004587I0000118J0000000D01*
G01X0001181Y0004351D02*
G03X0001299Y0004469I0000000J0000118D01*
G01X0001063D02*
G03X0001181Y0004351I0000118J0000000D01*
Y0004587D02*
G03X0001063Y0004469I0000000J0000118D01*
G01X0001299D02*
G03X0001181Y0004587I0000118J0000000D01*
G01X0012283Y0004351D02*
G03X0012401Y0004469I0000000J0000118D01*
G01X0012165D02*
G03X0012283Y0004351I0000118J0000000D01*
Y0004588D02*
G03X0012164Y0004469I0000000J0000119D01*
G01X0012402D02*
G03X0012283Y0004588I0000119J0000000D01*
G01X0001181Y-0006752D02*
G03X0001299Y-0006634I0000000J0000118D01*
G01X0001063D02*
G03X0001181Y-0006752I0000118J0000000D01*
Y-0006516D02*
G03X0001063Y-0006634I0000000J0000118D01*
G01X0001299D02*
G03X0001181Y-0006516I0000118J0000000D01*
G01X-0021024Y-0006752D02*
G03X-0020906Y-0006634I0000000J0000118D01*
G01X-0021142D02*
G03X-0021024Y-0006752I0000118J0000000D01*
Y-0006516D02*
G03X-0021142Y-0006634I0000000J0000118D01*
G01X-0020906D02*
G03X-0021024Y-0006516I0000118J0000000D01*
G01X-0009921Y-0006752D02*
G03X-0009803Y-0006634I0000000J0000118D01*
G01X-0010039D02*
G03X-0009921Y-0006752I0000118J0000000D01*
Y-0006516D02*
G03X-0010039Y-0006634I0000000J0000118D01*
G01X-0009803D02*
G03X-0009921Y-0006516I0000118J0000000D01*
G01X0012283Y-0006752D02*
G03X0012401Y-0006634I0000000J0000118D01*
G01X0012165D02*
G03X0012283Y-0006752I0000118J0000000D01*
Y-0006515D02*
G03X0012164Y-0006634I0000000J0000119D01*
G01X0012402D02*
G03X0012283Y-0006515I0000119J0000000D01*
G01X-0021024Y0015453D02*
G03X-0020906Y0015571I0000000J0000118D01*
G01X-0021142D02*
G03X-0021024Y0015453I0000118J0000000D01*
Y0015689D02*
G03X-0021142Y0015571I0000000J0000118D01*
G01X-0020906D02*
G03X-0021024Y0015689I0000118J0000000D01*
G01X-0009921Y0015453D02*
G03X-0009803Y0015571I0000000J0000118D01*
G01X-0010039D02*
G03X-0009921Y0015453I0000118J0000000D01*
Y0015689D02*
G03X-0010039Y0015571I0000000J0000118D01*
G01X-0009803D02*
G03X-0009921Y0015689I0000118J0000000D01*
G01X0001181Y0015453D02*
G03X0001299Y0015571I0000000J0000118D01*
G01X0001063D02*
G03X0001181Y0015453I0000118J0000000D01*
Y0015689D02*
G03X0001063Y0015571I0000000J0000118D01*
G01X0001299D02*
G03X0001181Y0015689I0000118J0000000D01*
G01X0012283Y0015453D02*
G03X0012401Y0015571I0000000J0000118D01*
G01X0012165D02*
G03X0012283Y0015453I0000118J0000000D01*
Y0015690D02*
G03X0012164Y0015571I0000000J0000119D01*
G01X0012402D02*
G03X0012283Y0015690I0000119J0000000D01*
G01X-0009921Y0026555D02*
G03X-0009803Y0026673I0000000J0000118D01*
G01X-0010039D02*
G03X-0009921Y0026555I0000118J0000000D01*
Y0026791D02*
G03X-0010039Y0026673I0000000J0000118D01*
G01X-0009803D02*
G03X-0009921Y0026791I0000118J0000000D01*
G01X-0021024Y0026555D02*
G03X-0020906Y0026673I0000000J0000118D01*
G01X-0021142D02*
G03X-0021024Y0026555I0000118J0000000D01*
Y0026791D02*
G03X-0021142Y0026673I0000000J0000118D01*
G01X-0020906D02*
G03X-0021024Y0026791I0000118J0000000D01*
G01X0001181Y0026555D02*
G03X0001299Y0026673I0000000J0000118D01*
G01X0001063D02*
G03X0001181Y0026555I0000118J0000000D01*
Y0026791D02*
G03X0001063Y0026673I0000000J0000118D01*
G01X0001299D02*
G03X0001181Y0026791I0000118J0000000D01*
G54D34*
G01X0018091Y0026997D02*
G03X0018141Y0027047I0000000J0000050D01*
G01X0018041D02*
G03X0018091Y0026997I0000050J0000000D01*
Y0027096D02*
G03X0018042Y0027047I0000000J0000049D01*
G01X0018140D02*
G03X0018091Y0027096I0000049J0000000D01*
G01X0015217Y0026997D02*
G03X0015267Y0027047I0000000J0000050D01*
G01X0015167D02*
G03X0015217Y0026997I0000050J0000000D01*
Y0027096D02*
G03X0015168Y0027047I0000000J0000049D01*
G01X0015266D02*
G03X0015217Y0027096I0000049J0000000D01*
G01X-0018091Y0004794D02*
G03X-0018042Y0004843I0000000J0000049D01*
G01X-0018140D02*
G03X-0018091Y0004794I0000049J0000000D01*
Y0004893D02*
G03X-0018141Y0004843I0000000J0000050D01*
G01X-0018041D02*
G03X-0018091Y0004893I0000050J0000000D01*
G01X-0015217Y0004794D02*
G03X-0015168Y0004843I0000000J0000049D01*
G01X-0015266D02*
G03X-0015217Y0004794I0000049J0000000D01*
Y0004893D02*
G03X-0015267Y0004843I0000000J0000050D01*
G01X-0015167D02*
G03X-0015217Y0004893I0000050J0000000D01*
G01X-0006988Y0004794D02*
G03X-0006939Y0004843I0000000J0000049D01*
G01X-0007037D02*
G03X-0006988Y0004794I0000049J0000000D01*
Y0004892D02*
G03X-0007037Y0004843I0000000J0000049D01*
G01X-0006939D02*
G03X-0006988Y0004892I0000049J0000000D01*
G01X-0004114Y0004794D02*
G03X-0004065Y0004843I0000000J0000049D01*
G01X-0004163D02*
G03X-0004114Y0004794I0000049J0000000D01*
Y0004892D02*
G03X-0004163Y0004843I0000000J0000049D01*
G01X-0004065D02*
G03X-0004114Y0004892I0000049J0000000D01*
G01X0004114Y0004794D02*
G03X0004163Y0004843I0000000J0000049D01*
G01X0004065D02*
G03X0004114Y0004794I0000049J0000000D01*
Y0004892D02*
G03X0004065Y0004843I0000000J0000049D01*
G01X0004163D02*
G03X0004114Y0004892I0000049J0000000D01*
G01X0006988Y0004794D02*
G03X0007037Y0004843I0000000J0000049D01*
G01X0006939D02*
G03X0006988Y0004794I0000049J0000000D01*
Y0004892D02*
G03X0006939Y0004843I0000000J0000049D01*
G01X0007037D02*
G03X0006988Y0004892I0000049J0000000D01*
G01X0015217Y0004793D02*
G03X0015267Y0004843I0000000J0000050D01*
G01X0015167D02*
G03X0015217Y0004793I0000050J0000000D01*
Y0004892D02*
G03X0015168Y0004843I0000000J0000049D01*
G01X0015266D02*
G03X0015217Y0004892I0000049J0000000D01*
G01X0018091Y0004793D02*
G03X0018141Y0004843I0000000J0000050D01*
G01X0018041D02*
G03X0018091Y0004793I0000050J0000000D01*
Y0004892D02*
G03X0018042Y0004843I0000000J0000049D01*
G01X0018140D02*
G03X0018091Y0004892I0000049J0000000D01*
G01X0004114Y-0006309D02*
G03X0004163Y-0006260I0000000J0000049D01*
G01X0004065D02*
G03X0004114Y-0006309I0000049J0000000D01*
Y-0006211D02*
G03X0004065Y-0006260I0000000J0000049D01*
G01X0004163D02*
G03X0004114Y-0006211I0000049J0000000D01*
G01X0006988Y-0006309D02*
G03X0007037Y-0006260I0000000J0000049D01*
G01X0006939D02*
G03X0006988Y-0006309I0000049J0000000D01*
Y-0006211D02*
G03X0006939Y-0006260I0000000J0000049D01*
G01X0007037D02*
G03X0006988Y-0006211I0000049J0000000D01*
G01X-0018091Y-0006309D02*
G03X-0018042Y-0006260I0000000J0000049D01*
G01X-0018140D02*
G03X-0018091Y-0006309I0000049J0000000D01*
Y-0006210D02*
G03X-0018141Y-0006260I0000000J0000050D01*
G01X-0018041D02*
G03X-0018091Y-0006210I0000050J0000000D01*
G01X-0015217Y-0006309D02*
G03X-0015168Y-0006260I0000000J0000049D01*
G01X-0015266D02*
G03X-0015217Y-0006309I0000049J0000000D01*
Y-0006210D02*
G03X-0015267Y-0006260I0000000J0000050D01*
G01X-0015167D02*
G03X-0015217Y-0006210I0000050J0000000D01*
G01X-0006988Y-0006309D02*
G03X-0006939Y-0006260I0000000J0000049D01*
G01X-0007037D02*
G03X-0006988Y-0006309I0000049J0000000D01*
Y-0006211D02*
G03X-0007037Y-0006260I0000000J0000049D01*
G01X-0006939D02*
G03X-0006988Y-0006211I0000049J0000000D01*
G01X-0004114Y-0006309D02*
G03X-0004065Y-0006260I0000000J0000049D01*
G01X-0004163D02*
G03X-0004114Y-0006309I0000049J0000000D01*
Y-0006211D02*
G03X-0004163Y-0006260I0000000J0000049D01*
G01X-0004065D02*
G03X-0004114Y-0006211I0000049J0000000D01*
G01X0015217Y-0006310D02*
G03X0015267Y-0006260I0000000J0000050D01*
G01X0015167D02*
G03X0015217Y-0006310I0000050J0000000D01*
Y-0006211D02*
G03X0015168Y-0006260I0000000J0000049D01*
G01X0015266D02*
G03X0015217Y-0006211I0000049J0000000D01*
G01X0018091Y-0006310D02*
G03X0018141Y-0006260I0000000J0000050D01*
G01X0018041D02*
G03X0018091Y-0006310I0000050J0000000D01*
Y-0006211D02*
G03X0018042Y-0006260I0000000J0000049D01*
G01X0018140D02*
G03X0018091Y-0006211I0000049J0000000D01*
G01X-0018091Y0015896D02*
G03X-0018042Y0015945I0000000J0000049D01*
G01X-0018140D02*
G03X-0018091Y0015896I0000049J0000000D01*
Y0015995D02*
G03X-0018141Y0015945I0000000J0000050D01*
G01X-0018041D02*
G03X-0018091Y0015995I0000050J0000000D01*
G01X-0015217Y0015896D02*
G03X-0015168Y0015945I0000000J0000049D01*
G01X-0015266D02*
G03X-0015217Y0015896I0000049J0000000D01*
Y0015995D02*
G03X-0015267Y0015945I0000000J0000050D01*
G01X-0015167D02*
G03X-0015217Y0015995I0000050J0000000D01*
G01X-0006988Y0015896D02*
G03X-0006939Y0015945I0000000J0000049D01*
G01X-0007037D02*
G03X-0006988Y0015896I0000049J0000000D01*
Y0015994D02*
G03X-0007037Y0015945I0000000J0000049D01*
G01X-0006939D02*
G03X-0006988Y0015994I0000049J0000000D01*
G01X-0004114Y0015896D02*
G03X-0004065Y0015945I0000000J0000049D01*
G01X-0004163D02*
G03X-0004114Y0015896I0000049J0000000D01*
Y0015994D02*
G03X-0004163Y0015945I0000000J0000049D01*
G01X-0004065D02*
G03X-0004114Y0015994I0000049J0000000D01*
G01X0004114Y0015896D02*
G03X0004163Y0015945I0000000J0000049D01*
G01X0004065D02*
G03X0004114Y0015896I0000049J0000000D01*
Y0015994D02*
G03X0004065Y0015945I0000000J0000049D01*
G01X0004163D02*
G03X0004114Y0015994I0000049J0000000D01*
G01X0006988Y0015896D02*
G03X0007037Y0015945I0000000J0000049D01*
G01X0006939D02*
G03X0006988Y0015896I0000049J0000000D01*
Y0015994D02*
G03X0006939Y0015945I0000000J0000049D01*
G01X0007037D02*
G03X0006988Y0015994I0000049J0000000D01*
G01X0015217Y0015895D02*
G03X0015267Y0015945I0000000J0000050D01*
G01X0015167D02*
G03X0015217Y0015895I0000050J0000000D01*
Y0015994D02*
G03X0015168Y0015945I0000000J0000049D01*
G01X0015266D02*
G03X0015217Y0015994I0000049J0000000D01*
G01X0018091Y0015895D02*
G03X0018141Y0015945I0000000J0000050D01*
G01X0018041D02*
G03X0018091Y0015895I0000050J0000000D01*
Y0015994D02*
G03X0018042Y0015945I0000000J0000049D01*
G01X0018140D02*
G03X0018091Y0015994I0000049J0000000D01*
G01X-0006988Y0026998D02*
G03X-0006939Y0027047I0000000J0000049D01*
G01X-0007037D02*
G03X-0006988Y0026998I0000049J0000000D01*
Y0027096D02*
G03X-0007037Y0027047I0000000J0000049D01*
G01X-0006939D02*
G03X-0006988Y0027096I0000049J0000000D01*
G01X-0004114Y0026998D02*
G03X-0004065Y0027047I0000000J0000049D01*
G01X-0004163D02*
G03X-0004114Y0026998I0000049J0000000D01*
Y0027096D02*
G03X-0004163Y0027047I0000000J0000049D01*
G01X-0004065D02*
G03X-0004114Y0027096I0000049J0000000D01*
G01X-0018091Y0026998D02*
G03X-0018042Y0027047I0000000J0000049D01*
G01X-0018140D02*
G03X-0018091Y0026998I0000049J0000000D01*
Y0027097D02*
G03X-0018141Y0027047I0000000J0000050D01*
G01X-0018041D02*
G03X-0018091Y0027097I0000050J0000000D01*
G01X-0015217Y0026998D02*
G03X-0015168Y0027047I0000000J0000049D01*
G01X-0015266D02*
G03X-0015217Y0026998I0000049J0000000D01*
Y0027097D02*
G03X-0015267Y0027047I0000000J0000050D01*
G01X-0015167D02*
G03X-0015217Y0027097I0000050J0000000D01*
G01X0006988Y0026998D02*
G03X0007037Y0027047I0000000J0000049D01*
G01X0006939D02*
G03X0006988Y0026998I0000049J0000000D01*
Y0027096D02*
G03X0006939Y0027047I0000000J0000049D01*
G01X0007037D02*
G03X0006988Y0027096I0000049J0000000D01*
G01X0004114Y0026998D02*
G03X0004163Y0027047I0000000J0000049D01*
G01X0004065D02*
G03X0004114Y0026998I0000049J0000000D01*
Y0027096D02*
G03X0004065Y0027047I0000000J0000049D01*
G01X0004163D02*
G03X0004114Y0027096I0000049J0000000D01*
G54D156*
G01X0017283Y-0018828D02*
Y-0019097D01*
X0017248Y-0018898D02*
Y-0019167D01*
X0017214Y-0018967D02*
Y-0019236D01*
X0017179Y-0019037D02*
Y-0019306D01*
X0017144Y-0019106D02*
Y-0019375D01*
X0017110Y-0019176D02*
Y-0019444D01*
X0017075Y-0019245D02*
Y-0019514D01*
X0017040Y-0019314D02*
Y-0019583D01*
X0017006Y-0019383D02*
Y-0019653D01*
X0016971Y-0019453D02*
Y-0019722D01*
X0016936Y-0019522D02*
Y-0019792D01*
X0016902Y-0019592D02*
Y-0019861D01*
X0016867Y-0019551D02*
Y-0019820D01*
X0016832Y-0019482D02*
Y-0019751D01*
X0016797Y-0019412D02*
Y-0019681D01*
X0016763Y-0019343D02*
Y-0019612D01*
X0016728Y-0019274D02*
Y-0019543D01*
X0016693Y-0019204D02*
Y-0019473D01*
X0016659Y-0019135D02*
Y-0019404D01*
X0016624Y-0019065D02*
Y-0019334D01*
X0016589Y-0018996D02*
Y-0019265D01*
X0016555Y-0018927D02*
Y-0019195D01*
X0016520Y-0018857D02*
Y-0019126D01*
X0016485Y-0018788D02*
Y-0019140D01*
X0016450Y-0018719D02*
Y-0019554D01*
X0016416Y-0018649D02*
Y-0019876D01*
X0016381Y-0018580D02*
Y-0019876D01*
X0016346Y-0018632D02*
Y-0019876D01*
X0016312Y-0018978D02*
Y-0019876D01*
X0016277Y-0019325D02*
Y-0019876D01*
X0016242Y-0019671D02*
Y-0019876D01*
X0016377Y-0018571D02*
X0016352D01*
X0016394Y-0018606D02*
X0016349D01*
X0016411Y-0018641D02*
X0016345D01*
X0016429Y-0018675D02*
X0016342D01*
X0016446Y-0018710D02*
X0016339D01*
X0016464Y-0018745D02*
X0016335D01*
X0016481Y-0018780D02*
X0016331D01*
X0016498Y-0018814D02*
X0016328D01*
X0016516Y-0018849D02*
X0016325D01*
X0016533Y-0018883D02*
X0016321D01*
X0016550Y-0018918D02*
X0016318D01*
X0016568Y-0018953D02*
X0016314D01*
X0016585Y-0018988D02*
X0016311D01*
X0016602Y-0019022D02*
X0016307D01*
X0016620Y-0019057D02*
X0016304D01*
X0016489Y-0019092D02*
X0016300D01*
X0016486Y-0019126D02*
X0016297D01*
X0016483Y-0019161D02*
X0016293D01*
X0016480Y-0019196D02*
X0016290D01*
X0016478Y-0019230D02*
X0016287D01*
X0016475Y-0019265D02*
X0016283D01*
X0016472Y-0019300D02*
X0016280D01*
X0016469Y-0019335D02*
X0016276D01*
X0016466Y-0019369D02*
X0016272D01*
X0016463Y-0019404D02*
X0016269D01*
X0016460Y-0019439D02*
X0016266D01*
X0016457Y-0019473D02*
X0016262D01*
X0016454Y-0019508D02*
X0016259D01*
X0016451Y-0019543D02*
X0016255D01*
X0016448Y-0019578D02*
X0016252D01*
X0016446Y-0019612D02*
X0016248D01*
X0016443Y-0019647D02*
X0016245D01*
X0016440Y-0019681D02*
X0016241D01*
X0016437Y-0019716D02*
X0016238D01*
X0016434Y-0019751D02*
X0016234D01*
X0016431Y-0019785D02*
X0016231D01*
X0016428Y-0019820D02*
X0016228D01*
X0017502Y-0019230D02*
X0017311D01*
X0017217D02*
X0017082D01*
X0016706D02*
X0016572D01*
X0017506Y-0019265D02*
X0017314D01*
X0017199D02*
X0017065D01*
X0016724D02*
X0016589D01*
X0017509Y-0019300D02*
X0017317D01*
X0017182D02*
X0017047D01*
X0016741D02*
X0016607D01*
X0017513Y-0019335D02*
X0017320D01*
X0017165D02*
X0017030D01*
X0016759D02*
X0016624D01*
X0017516Y-0019369D02*
X0017323D01*
X0017147D02*
X0017013D01*
X0016776D02*
X0016641D01*
X0017520Y-0019404D02*
X0017326D01*
X0017130D02*
X0016995D01*
X0016793D02*
X0016659D01*
X0017523Y-0019439D02*
X0017328D01*
X0017113D02*
X0016978D01*
X0016811D02*
X0016676D01*
X0017526Y-0019473D02*
X0017331D01*
X0017095D02*
X0016961D01*
X0016828D02*
X0016693D01*
X0017530Y-0019508D02*
X0017334D01*
X0017078D02*
X0016943D01*
X0016845D02*
X0016711D01*
X0017533Y-0019543D02*
X0017337D01*
X0017061D02*
X0016926D01*
X0016863D02*
X0016728D01*
X0017537Y-0019578D02*
X0017340D01*
X0017043D02*
X0016909D01*
X0016880D02*
X0016745D01*
X0017541Y-0019612D02*
X0017343D01*
X0017026D02*
X0016763D01*
X0017544Y-0019647D02*
X0017346D01*
X0017009D02*
X0016780D01*
X0017547Y-0019681D02*
X0017349D01*
X0016991D02*
X0016797D01*
X0017551Y-0019716D02*
X0017352D01*
X0016974D02*
X0016815D01*
X0017554Y-0019751D02*
X0017355D01*
X0016956D02*
X0016832D01*
X0017558Y-0019785D02*
X0017357D01*
X0016939D02*
X0016850D01*
X0017561Y-0019820D02*
X0017361D01*
X0016922D02*
X0016867D01*
X0017565Y-0019855D02*
X0017363D01*
X0016904D02*
X0016884D01*
X0016425D02*
X0016224D01*
X0016424Y-0019876D02*
X0016222D01*
X0016491Y-0019069D02*
X0016424Y-0019876D01*
X0016491Y-0019069D02*
X0016894Y-0019876D01*
X0017298Y-0019069D02*
X0016894Y-0019876D01*
X0017298Y-0019069D02*
X0017365Y-0019876D01*
X0017567D02*
X0017365D01*
X0017432Y-0018531D02*
X0017567Y-0019876D01*
X0017432Y-0018531D02*
X0016894Y-0019606D01*
X0016357Y-0018531D02*
X0016894Y-0019606D01*
X0016357Y-0018531D02*
X0016222Y-0019876D01*
X0017561Y-0019815D02*
Y-0019876D01*
X0017526Y-0019469D02*
Y-0019876D01*
X0017491Y-0019122D02*
Y-0019876D01*
X0017457Y-0018775D02*
Y-0019876D01*
X0017422Y-0018551D02*
Y-0019876D01*
X0017387Y-0018620D02*
Y-0019876D01*
X0017352Y-0018690D02*
Y-0019725D01*
X0017318Y-0018759D02*
Y-0019311D01*
X0017436Y-0018571D02*
X0017412D01*
X0017440Y-0018606D02*
X0017394D01*
X0017443Y-0018641D02*
X0017377D01*
X0017446Y-0018675D02*
X0017360D01*
X0017450Y-0018710D02*
X0017343D01*
X0017454Y-0018745D02*
X0017325D01*
X0017457Y-0018780D02*
X0017307D01*
X0017461Y-0018814D02*
X0017290D01*
X0017464Y-0018849D02*
X0017273D01*
X0017467Y-0018883D02*
X0017256D01*
X0017471Y-0018918D02*
X0017238D01*
X0017474Y-0018953D02*
X0017221D01*
X0017478Y-0018988D02*
X0017204D01*
X0017481Y-0019022D02*
X0017186D01*
X0017485Y-0019057D02*
X0017169D01*
X0017488Y-0019092D02*
X0017299D01*
X0017286D02*
X0017152D01*
X0016637D02*
X0016503D01*
X0017492Y-0019126D02*
X0017302D01*
X0017269D02*
X0017134D01*
X0016654D02*
X0016520D01*
X0017495Y-0019161D02*
X0017305D01*
X0017251D02*
X0017117D01*
X0016672D02*
X0016537D01*
X0017499Y-0019196D02*
X0017308D01*
X0017234D02*
X0017100D01*
X0016689D02*
X0016555D01*
X0015522Y-0018531D02*
Y-0019876D01*
X0015487Y-0018531D02*
Y-0019876D01*
X0015452Y-0018531D02*
Y-0019876D01*
X0015418Y-0018531D02*
Y-0019876D01*
X0015383Y-0018531D02*
Y-0019876D01*
X0015348Y-0018531D02*
Y-0019876D01*
X0015314Y-0018531D02*
Y-0019876D01*
X0015279Y-0018531D02*
Y-0018800D01*
X0015244Y-0018531D02*
Y-0018800D01*
X0015210Y-0018531D02*
Y-0018800D01*
X0015175Y-0018531D02*
Y-0018800D01*
X0015140Y-0018531D02*
Y-0018800D01*
X0015106Y-0018531D02*
Y-0018800D01*
X0015071Y-0018531D02*
Y-0018800D01*
X0015036Y-0018531D02*
Y-0018800D01*
X0015002Y-0018531D02*
Y-0018800D01*
X0014967Y-0018531D02*
Y-0018800D01*
X0014932Y-0018531D02*
Y-0018800D01*
X0014897Y-0018531D02*
Y-0018800D01*
X0015953Y-0018537D02*
X0014877D01*
X0015953Y-0018571D02*
X0014877D01*
X0015953Y-0018606D02*
X0014877D01*
X0015953Y-0018641D02*
X0014877D01*
X0015953Y-0018675D02*
X0014877D01*
X0015953Y-0018710D02*
X0014877D01*
X0015953Y-0018745D02*
X0014877D01*
X0015953Y-0018780D02*
X0014877D01*
X0015550Y-0018814D02*
X0015280D01*
X0015550Y-0018849D02*
X0015280D01*
X0015550Y-0018883D02*
X0015280D01*
X0015550Y-0018918D02*
X0015280D01*
X0015550Y-0018953D02*
X0015280D01*
X0015550Y-0018988D02*
X0015280D01*
X0015550Y-0019022D02*
X0015280D01*
X0015550Y-0019057D02*
X0015280D01*
X0015550Y-0019092D02*
X0015280D01*
X0015550Y-0019126D02*
X0015280D01*
X0015550Y-0019161D02*
X0015280D01*
X0015550Y-0019196D02*
X0015280D01*
X0015550Y-0019230D02*
X0015280D01*
X0015550Y-0019265D02*
X0015280D01*
X0015550Y-0019300D02*
X0015280D01*
X0015550Y-0019335D02*
X0015280D01*
X0015550Y-0019369D02*
X0015280D01*
X0015550Y-0019404D02*
X0015280D01*
X0015550Y-0019439D02*
X0015280D01*
X0015550Y-0019473D02*
X0015280D01*
X0015550Y-0019508D02*
X0015280D01*
X0015550Y-0019543D02*
X0015280D01*
X0015550Y-0019578D02*
X0015280D01*
X0015550Y-0019612D02*
X0015280D01*
X0015550Y-0019647D02*
X0015280D01*
X0015550Y-0019681D02*
X0015280D01*
X0015550Y-0019716D02*
X0015280D01*
X0015550Y-0019751D02*
X0015280D01*
X0015550Y-0019785D02*
X0015280D01*
X0015550Y-0019820D02*
X0015280D01*
X0015550Y-0019855D02*
X0015280D01*
X0015953Y-0018531D02*
X0014877D01*
X0015953D02*
Y-0018800D01*
X0015550D01*
Y-0019876D01*
X0015280D01*
Y-0018800D02*
Y-0019876D01*
Y-0018800D02*
X0014877D01*
Y-0018531D02*
Y-0018800D01*
X0015938Y-0018531D02*
Y-0018800D01*
X0015904Y-0018531D02*
Y-0018800D01*
X0015869Y-0018531D02*
Y-0018800D01*
X0015834Y-0018531D02*
Y-0018800D01*
X0015800Y-0018531D02*
Y-0018800D01*
X0015765Y-0018531D02*
Y-0018800D01*
X0015730Y-0018531D02*
Y-0018800D01*
X0015695Y-0018531D02*
Y-0018800D01*
X0015661Y-0018531D02*
Y-0018800D01*
X0015626Y-0018531D02*
Y-0018800D01*
X0015591Y-0018531D02*
Y-0018800D01*
X0015557Y-0018531D02*
Y-0018800D01*
X0013253Y-0019548D02*
Y-0020696D01*
Y-0023177D02*
Y-0024845D01*
X0013218Y-0019520D02*
Y-0020719D01*
Y-0023156D02*
Y-0024640D01*
X0013183Y-0019491D02*
Y-0020740D01*
Y-0023134D02*
Y-0024499D01*
X0013149Y-0019463D02*
Y-0020736D01*
Y-0023113D02*
Y-0024431D01*
X0013114Y-0019435D02*
Y-0020682D01*
Y-0023092D02*
Y-0024363D01*
X0013080Y-0019414D02*
Y-0020628D01*
Y-0023070D02*
Y-0024295D01*
X0013044Y-0019395D02*
Y-0020573D01*
Y-0023049D02*
Y-0024227D01*
X0013010Y-0019376D02*
Y-0020519D01*
Y-0023028D02*
Y-0024182D01*
X0012975Y-0019357D02*
Y-0020474D01*
Y-0023006D02*
Y-0024144D01*
X0012941Y-0019338D02*
Y-0020433D01*
Y-0022985D02*
Y-0024107D01*
X0012906Y-0019319D02*
Y-0020391D01*
Y-0022964D02*
Y-0024070D01*
X0012871Y-0019300D02*
Y-0020350D01*
Y-0022943D02*
Y-0024033D01*
X0012837Y-0019281D02*
Y-0020309D01*
Y-0022922D02*
Y-0023995D01*
X0012802Y-0019262D02*
Y-0020274D01*
Y-0022905D02*
Y-0023958D01*
X0012767Y-0019243D02*
Y-0020244D01*
Y-0022888D02*
Y-0023931D01*
X0012732Y-0019228D02*
Y-0020215D01*
Y-0022871D02*
Y-0023906D01*
X0012698Y-0019217D02*
Y-0020185D01*
Y-0022854D02*
Y-0023882D01*
X0012663Y-0019205D02*
Y-0020155D01*
Y-0022837D02*
Y-0023857D01*
X0012628Y-0019193D02*
Y-0020126D01*
Y-0022820D02*
Y-0023832D01*
X0012594Y-0019181D02*
Y-0020104D01*
Y-0022803D02*
Y-0023807D01*
X0012559Y-0019170D02*
Y-0020085D01*
Y-0022786D02*
Y-0023783D01*
X0012524Y-0019158D02*
Y-0020065D01*
Y-0022769D02*
Y-0023758D01*
X0012489Y-0019146D02*
Y-0020046D01*
Y-0022752D02*
Y-0023735D01*
X0012455Y-0019135D02*
Y-0020027D01*
Y-0022735D02*
Y-0023717D01*
X0012420Y-0019123D02*
Y-0020007D01*
Y-0022718D02*
Y-0023698D01*
X0012385Y-0019111D02*
Y-0019990D01*
Y-0022701D02*
Y-0023680D01*
X0012351Y-0019103D02*
Y-0019979D01*
Y-0022685D02*
Y-0023661D01*
X0012316Y-0019098D02*
Y-0019968D01*
Y-0022669D02*
Y-0023642D01*
X0012281Y-0019093D02*
Y-0019957D01*
Y-0022654D02*
Y-0023624D01*
X0012247Y-0019088D02*
Y-0019946D01*
Y-0022639D02*
Y-0023605D01*
X0012212Y-0019083D02*
Y-0019935D01*
Y-0022623D02*
Y-0023587D01*
X0012177Y-0019078D02*
Y-0019924D01*
Y-0022608D02*
Y-0023568D01*
X0012143Y-0019072D02*
Y-0019913D01*
Y-0022592D02*
Y-0023551D01*
X0012108Y-0019067D02*
Y-0019907D01*
Y-0022577D02*
Y-0023535D01*
X0012073Y-0019062D02*
Y-0019904D01*
Y-0022561D02*
Y-0023518D01*
X0012039Y-0019057D02*
Y-0019900D01*
Y-0022546D02*
Y-0023502D01*
X0012004Y-0019052D02*
Y-0019896D01*
Y-0022531D02*
Y-0023486D01*
X0011969Y-0019047D02*
Y-0019892D01*
Y-0022515D02*
Y-0023469D01*
X0011934Y-0019044D02*
Y-0019888D01*
Y-0022500D02*
Y-0023453D01*
X0011900Y-0019046D02*
Y-0019884D01*
Y-0022484D02*
Y-0023437D01*
X0011865Y-0019047D02*
Y-0019880D01*
Y-0022469D02*
Y-0023420D01*
X0011830Y-0019048D02*
Y-0019876D01*
Y-0022454D02*
Y-0023404D01*
X0011796Y-0019050D02*
Y-0019879D01*
Y-0022439D02*
Y-0023388D01*
X0011761Y-0019051D02*
Y-0019881D01*
Y-0022424D02*
Y-0023374D01*
X0011726Y-0019052D02*
Y-0019884D01*
Y-0022409D02*
Y-0023359D01*
X0011692Y-0019053D02*
Y-0019886D01*
Y-0022393D02*
Y-0023343D01*
X0011657Y-0019055D02*
Y-0019889D01*
Y-0022378D02*
Y-0023328D01*
X0011622Y-0019056D02*
Y-0019892D01*
Y-0022362D02*
Y-0023313D01*
X0011587Y-0019057D02*
Y-0019894D01*
Y-0022346D02*
Y-0023298D01*
X0011553Y-0019058D02*
Y-0019897D01*
Y-0022331D02*
Y-0023282D01*
X0011518Y-0019059D02*
Y-0019899D01*
Y-0022314D02*
Y-0023267D01*
X0011483Y-0019061D02*
Y-0019904D01*
Y-0022297D02*
Y-0023252D01*
X0011449Y-0019062D02*
Y-0019915D01*
Y-0022280D02*
Y-0023237D01*
X0011414Y-0019067D02*
Y-0019925D01*
Y-0022263D02*
Y-0023222D01*
X0011379Y-0019076D02*
Y-0019936D01*
Y-0022246D02*
Y-0023207D01*
X0011344Y-0019084D02*
Y-0019947D01*
Y-0022230D02*
Y-0023192D01*
X0011310Y-0019093D02*
Y-0019958D01*
Y-0022213D02*
Y-0023177D01*
X0011275Y-0019102D02*
Y-0019969D01*
Y-0022196D02*
Y-0023162D01*
X0011241Y-0019110D02*
Y-0019980D01*
Y-0022177D02*
Y-0023145D01*
X0011206Y-0019119D02*
Y-0019991D01*
Y-0022156D02*
Y-0023129D01*
X0011171Y-0019128D02*
Y-0020003D01*
Y-0022136D02*
Y-0023113D01*
X0011137Y-0019136D02*
Y-0020024D01*
Y-0022115D02*
Y-0023096D01*
X0011102Y-0019145D02*
Y-0020044D01*
Y-0022095D02*
Y-0023080D01*
X0011067Y-0019154D02*
Y-0020065D01*
Y-0022075D02*
Y-0023063D01*
X0011032Y-0019162D02*
Y-0020086D01*
Y-0022054D02*
Y-0023046D01*
X0010998Y-0019171D02*
Y-0020107D01*
Y-0022034D02*
Y-0023030D01*
X0010963Y-0019180D02*
Y-0020128D01*
Y-0022008D02*
Y-0023014D01*
X0010928Y-0019188D02*
Y-0020148D01*
Y-0021980D02*
Y-0022996D01*
X0010894Y-0019197D02*
Y-0020170D01*
Y-0021953D02*
Y-0022976D01*
X0010859Y-0019213D02*
Y-0020206D01*
Y-0021925D02*
Y-0022957D01*
X0010824Y-0019231D02*
Y-0020241D01*
Y-0021897D02*
Y-0022938D01*
X0010789Y-0019249D02*
Y-0020276D01*
Y-0021869D02*
Y-0022919D01*
X0010755Y-0019267D02*
Y-0020310D01*
Y-0021842D02*
Y-0022899D01*
X0010720Y-0019285D02*
Y-0020345D01*
Y-0021802D02*
Y-0022880D01*
X0010685Y-0019302D02*
Y-0020380D01*
Y-0021760D02*
Y-0022861D01*
X0010651Y-0019320D02*
Y-0020431D01*
Y-0021717D02*
Y-0022842D01*
X0010616Y-0019338D02*
Y-0020492D01*
Y-0021675D02*
Y-0022822D01*
X0010581Y-0019356D02*
Y-0020553D01*
Y-0021633D02*
Y-0022803D01*
X0010546Y-0019374D02*
Y-0020614D01*
Y-0021573D02*
Y-0022784D01*
X0010512Y-0019391D02*
Y-0020678D01*
Y-0021486D02*
Y-0022761D01*
X0010477Y-0019409D02*
Y-0020821D01*
Y-0021399D02*
Y-0022736D01*
X0010443Y-0019427D02*
Y-0020964D01*
Y-0021176D02*
Y-0022711D01*
X0010408Y-0019444D02*
Y-0022686D01*
X0010373Y-0019474D02*
Y-0022661D01*
X0010339Y-0019505D02*
Y-0022635D01*
X0010304Y-0019535D02*
Y-0022610D01*
X0010269Y-0019565D02*
Y-0022585D01*
X0010234Y-0019596D02*
Y-0022560D01*
X0010200Y-0019626D02*
Y-0022535D01*
X0010165Y-0019657D02*
Y-0022509D01*
X0010130Y-0019687D02*
Y-0022473D01*
X0010096Y-0019717D02*
Y-0022436D01*
X0010061Y-0019748D02*
Y-0022399D01*
X0010026Y-0019778D02*
Y-0022362D01*
X0009991Y-0019819D02*
Y-0022324D01*
X0009957Y-0019871D02*
Y-0022287D01*
X0009922Y-0019924D02*
Y-0022250D01*
X0009887Y-0019977D02*
Y-0022213D01*
X0009853Y-0020030D02*
Y-0022168D01*
X0009818Y-0020082D02*
Y-0022105D01*
X0009783Y-0020135D02*
Y-0022043D01*
X0009749Y-0020188D02*
Y-0021980D01*
X0009714Y-0020244D02*
Y-0021917D01*
X0009679Y-0020356D02*
Y-0021855D01*
X0009644Y-0020468D02*
Y-0021778D01*
X0009610Y-0020581D02*
Y-0021633D01*
X0009575Y-0020693D02*
Y-0021487D01*
X0009541Y-0021250D02*
Y-0021342D01*
X0013595Y-0019885D02*
X0011903D01*
X0013625Y-0019919D02*
X0012161D01*
X0013656Y-0019954D02*
X0012271D01*
X0013686Y-0019989D02*
X0012382D01*
X0013710Y-0020023D02*
X0012449D01*
X0013731Y-0020058D02*
X0012511D01*
X0013753Y-0020093D02*
X0012573D01*
X0013774Y-0020128D02*
X0012630D01*
X0013796Y-0020162D02*
X0012671D01*
X0013817Y-0020197D02*
X0012711D01*
X0013839Y-0020231D02*
X0012752D01*
X0013860Y-0020266D02*
X0012793D01*
X0013868Y-0020301D02*
X0012830D01*
X0013814Y-0020335D02*
X0012859D01*
X0013759Y-0020370D02*
X0012888D01*
X0013704Y-0020405D02*
X0012917D01*
X0013650Y-0020440D02*
X0012946D01*
X0013596Y-0020474D02*
X0012976D01*
X0013543Y-0020509D02*
X0013004D01*
X0013489Y-0020544D02*
X0013026D01*
X0013435Y-0020578D02*
X0013048D01*
X0013381Y-0020613D02*
X0013070D01*
X0013327Y-0020648D02*
X0013092D01*
X0013273Y-0020683D02*
X0013115D01*
X0013220Y-0020717D02*
X0013137D01*
X0014147Y-0025089D02*
X0013251D01*
X0014142Y-0025124D02*
X0013247D01*
X0014137Y-0025158D02*
X0013244D01*
X0014132Y-0025193D02*
X0013240D01*
X0014127Y-0025228D02*
X0013237D01*
X0014122Y-0025262D02*
X0013233D01*
X0014117Y-0025297D02*
X0013229D01*
X0014111Y-0025331D02*
X0013226D01*
X0014106Y-0025366D02*
X0013220D01*
X0014101Y-0025401D02*
X0013206D01*
X0014096Y-0025436D02*
X0013192D01*
X0014091Y-0025470D02*
X0013178D01*
X0014086Y-0025505D02*
X0013164D01*
X0014081Y-0025540D02*
X0013150D01*
X0014076Y-0025574D02*
X0013136D01*
X0014068Y-0025609D02*
X0013122D01*
X0014053Y-0025644D02*
X0013108D01*
X0014038Y-0025679D02*
X0013094D01*
X0014023Y-0025713D02*
X0013080D01*
X0014008Y-0025748D02*
X0013062D01*
X0013993Y-0025783D02*
X0013035D01*
X0013978Y-0025817D02*
X0013009D01*
X0013963Y-0025852D02*
X0012983D01*
X0013948Y-0025887D02*
X0012956D01*
X0013933Y-0025921D02*
X0012930D01*
X0013918Y-0025956D02*
X0012903D01*
X0013903Y-0025991D02*
X0012877D01*
X0013888Y-0026026D02*
X0012850D01*
X0013873Y-0026060D02*
X0012822D01*
X0013858Y-0026095D02*
X0012778D01*
X0013843Y-0026130D02*
X0012735D01*
X0013828Y-0026164D02*
X0012691D01*
X0013806Y-0026199D02*
X0012648D01*
X0013779Y-0026234D02*
X0012604D01*
X0013752Y-0026269D02*
X0012560D01*
X0013725Y-0026303D02*
X0012517D01*
X0013698Y-0026338D02*
X0012446D01*
X0013670Y-0026372D02*
X0012371D01*
X0013643Y-0026407D02*
X0012296D01*
X0013616Y-0026442D02*
X0012222D01*
X0013589Y-0026476D02*
X0012147D01*
X0013562Y-0026511D02*
X0011979D01*
X0013535Y-0026546D02*
X0011806D01*
X0011844Y-0027379D02*
X0011447D01*
X0012999Y-0020502D02*
X0013161Y-0020754D01*
X0012821Y-0020291D02*
X0012999Y-0020502D01*
X0012621Y-0020120D02*
X0012821Y-0020291D01*
X0012393Y-0019992D02*
X0012621Y-0020120D01*
X0012131Y-0019910D02*
X0012393Y-0019992D01*
X0011829Y-0019876D02*
X0012131Y-0019910D01*
X0011829Y-0019876D02*
X0011491Y-0019902D01*
X0011175Y-0020001D01*
X0010898Y-0020167D01*
X0010672Y-0020394D01*
X0010513Y-0020672D01*
X0010435Y-0020998D01*
X0010450Y-0021329D01*
X0010560Y-0021606D01*
X0010748Y-0021836D01*
X0010988Y-0022028D01*
X0011260Y-0022188D01*
X0011540Y-0022325D01*
X0011701Y-0022398D01*
X0011766Y-0022426D01*
X0011876Y-0022474D01*
X0012006Y-0022531D01*
X0012124Y-0022584D01*
X0012207Y-0022621D01*
X0012355Y-0022687D01*
X0012840Y-0022924D01*
X0013276Y-0023191D01*
X0013646Y-0023511D01*
X0013930Y-0023897D01*
X0014110Y-0024369D01*
X0014169Y-0024946D01*
X0014072Y-0025598D01*
X0013822Y-0026180D01*
X0013439Y-0026669D01*
X0012945Y-0027047D01*
X0012362Y-0027298D01*
X0011713Y-0027399D01*
X0011098Y-0027352D02*
X0011713Y-0027399D01*
X0010552Y-0027182D02*
X0011098Y-0027352D01*
X0010074Y-0026902D02*
X0010552Y-0027182D01*
X0009674Y-0026520D02*
X0010074Y-0026902D01*
X0009365Y-0026048D02*
X0009674Y-0026520D01*
X0009154Y-0025498D02*
X0009365Y-0026048D01*
X0009139Y-0025302D02*
X0009154Y-0025498D01*
X0009269Y-0025265D02*
X0009139Y-0025302D01*
X0009462Y-0025211D02*
X0009269Y-0025265D01*
X0009673Y-0025152D02*
X0009462Y-0025211D01*
X0009858Y-0025100D02*
X0009673Y-0025152D01*
X0009972Y-0025069D02*
X0009858Y-0025100D01*
X0009972Y-0025069D02*
X0010027Y-0025261D01*
X0010161Y-0025630D01*
X0010365Y-0025956D01*
X0010631Y-0026226D01*
X0010955Y-0026424D01*
X0011327Y-0026539D01*
X0011738Y-0026560D01*
X0012143Y-0026479D02*
X0011738Y-0026560D01*
X0012511Y-0026308D02*
X0012143Y-0026479D01*
X0012827Y-0026057D02*
X0012511Y-0026308D01*
X0013070Y-0025738D02*
X0012827Y-0026057D01*
X0013223Y-0025359D02*
X0013070Y-0025738D01*
X0013268Y-0024932D02*
X0013223Y-0025359D01*
X0013200Y-0024531D02*
X0013268Y-0024932D01*
X0013036Y-0024210D02*
X0013200Y-0024531D01*
X0012796Y-0023952D02*
X0013036Y-0024210D01*
X0012499Y-0023740D02*
X0012796Y-0023952D01*
X0012160Y-0023559D02*
X0012499Y-0023740D01*
X0011801Y-0023391D02*
X0012160Y-0023559D01*
X0011747Y-0023368D02*
X0011801Y-0023391D01*
X0011664Y-0023331D02*
X0011747Y-0023368D01*
X0011550Y-0023281D02*
X0011664Y-0023331D01*
X0011434Y-0023231D02*
X0011550Y-0023281D01*
X0011338Y-0023189D02*
X0011434Y-0023231D01*
X0011287Y-0023168D02*
X0011338Y-0023189D01*
X0010949Y-0023007D02*
X0011287Y-0023168D01*
X0010531Y-0022776D02*
X0010949Y-0023007D01*
X0010164Y-0022509D02*
X0010531Y-0022776D01*
X0009865Y-0022189D02*
X0010164Y-0022509D01*
X0009650Y-0021802D02*
X0009865Y-0022189D01*
X0009539Y-0021333D02*
X0009650Y-0021802D01*
X0009553Y-0020766D02*
X0009539Y-0021333D01*
X0009716Y-0020239D02*
X0009553Y-0020766D01*
X0010007Y-0019795D02*
X0009716Y-0020239D01*
X0010406Y-0019446D02*
X0010007Y-0019795D01*
X0010889Y-0019198D02*
X0010406Y-0019446D01*
X0011431Y-0019063D02*
X0010889Y-0019198D01*
X0011950Y-0019044D02*
X0011431Y-0019063D01*
X0011950Y-0019044D02*
X0012367Y-0019106D01*
X0012754Y-0019235D01*
X0013107Y-0019429D01*
X0013421Y-0019685D01*
X0013694Y-0019998D01*
X0013878Y-0020294D01*
X0013811Y-0020338D01*
X0013674Y-0020424D01*
X0013504Y-0020535D01*
X0013338Y-0020641D01*
X0013212Y-0020723D01*
X0013161Y-0020754D01*
X0014155Y-0024812D02*
Y-0025037D01*
X0014120Y-0024469D02*
Y-0025272D01*
X0014085Y-0024304D02*
Y-0025508D01*
X0014051Y-0024213D02*
Y-0025648D01*
X0014016Y-0024122D02*
Y-0025728D01*
X0013981Y-0024032D02*
Y-0025809D01*
X0013947Y-0023941D02*
Y-0025890D01*
X0013912Y-0023872D02*
Y-0025970D01*
X0013877Y-0023826D02*
Y-0026051D01*
X0013843Y-0023778D02*
Y-0026131D01*
X0013808Y-0023731D02*
Y-0026197D01*
X0013773Y-0023684D02*
Y-0026241D01*
X0013739Y-0023637D02*
Y-0026286D01*
X0013704Y-0023590D02*
Y-0026330D01*
X0013669Y-0023543D02*
Y-0026374D01*
X0013635Y-0023501D02*
Y-0026419D01*
X0013600Y-0023471D02*
Y-0026463D01*
X0013565Y-0023441D02*
Y-0026507D01*
X0013530Y-0023411D02*
Y-0026552D01*
X0013496Y-0023381D02*
Y-0026596D01*
X0013461Y-0023351D02*
Y-0026640D01*
X0013426Y-0023321D02*
Y-0026678D01*
X0013392Y-0023291D02*
Y-0026705D01*
X0013357Y-0023261D02*
Y-0026731D01*
X0013322Y-0023231D02*
Y-0026758D01*
X0013287Y-0023201D02*
Y-0026785D01*
X0013253Y-0025072D02*
Y-0026811D01*
X0013218Y-0025370D02*
Y-0026838D01*
X0013183Y-0025456D02*
Y-0026864D01*
X0013149Y-0025542D02*
Y-0026891D01*
X0013114Y-0025628D02*
Y-0026917D01*
X0013080Y-0025714D02*
Y-0026944D01*
X0013044Y-0025771D02*
Y-0026970D01*
X0013010Y-0025816D02*
Y-0026997D01*
X0012975Y-0025862D02*
Y-0027024D01*
X0012941Y-0025907D02*
Y-0027049D01*
X0012906Y-0025953D02*
Y-0027064D01*
X0012871Y-0025998D02*
Y-0027079D01*
X0012837Y-0026044D02*
Y-0027094D01*
X0012802Y-0026076D02*
Y-0027108D01*
X0012767Y-0026104D02*
Y-0027123D01*
X0012732Y-0026131D02*
Y-0027138D01*
X0012698Y-0026159D02*
Y-0027153D01*
X0012663Y-0026187D02*
Y-0027168D01*
X0012628Y-0026214D02*
Y-0027183D01*
X0012594Y-0026242D02*
Y-0027198D01*
X0012559Y-0026269D02*
Y-0027213D01*
X0012524Y-0026297D02*
Y-0027228D01*
X0012489Y-0026318D02*
Y-0027243D01*
X0012455Y-0026333D02*
Y-0027257D01*
X0012420Y-0026350D02*
Y-0027272D01*
X0012385Y-0026366D02*
Y-0027287D01*
X0012351Y-0026382D02*
Y-0027299D01*
X0012316Y-0026398D02*
Y-0027305D01*
X0012281Y-0026414D02*
Y-0027310D01*
X0012247Y-0026430D02*
Y-0027315D01*
X0012212Y-0026446D02*
Y-0027321D01*
X0012177Y-0026462D02*
Y-0027326D01*
X0012143Y-0026478D02*
Y-0027332D01*
X0012108Y-0026485D02*
Y-0027337D01*
X0012073Y-0026493D02*
Y-0027343D01*
X0012039Y-0026499D02*
Y-0027348D01*
X0012004Y-0026506D02*
Y-0027354D01*
X0011969Y-0026513D02*
Y-0027359D01*
X0011934Y-0026520D02*
Y-0027365D01*
X0011900Y-0026527D02*
Y-0027370D01*
X0011865Y-0026534D02*
Y-0027375D01*
X0011830Y-0026541D02*
Y-0027381D01*
X0011796Y-0026548D02*
Y-0027386D01*
X0011761Y-0026555D02*
Y-0027392D01*
X0011726Y-0026559D02*
Y-0027397D01*
X0011692Y-0026557D02*
Y-0027397D01*
X0011657Y-0026556D02*
Y-0027395D01*
X0011622Y-0026554D02*
Y-0027392D01*
X0011587Y-0026552D02*
Y-0027389D01*
X0011553Y-0026550D02*
Y-0027387D01*
X0011518Y-0026549D02*
Y-0027384D01*
X0011483Y-0026547D02*
Y-0027381D01*
X0011449Y-0026545D02*
Y-0027379D01*
X0011414Y-0026544D02*
Y-0027376D01*
X0011379Y-0026542D02*
Y-0027373D01*
X0011344Y-0026540D02*
Y-0027371D01*
X0011310Y-0026534D02*
Y-0027368D01*
X0011275Y-0026523D02*
Y-0027365D01*
X0011241Y-0026513D02*
Y-0027363D01*
X0011206Y-0026502D02*
Y-0027360D01*
X0011171Y-0026491D02*
Y-0027357D01*
X0011137Y-0026480D02*
Y-0027355D01*
X0011102Y-0026470D02*
Y-0027352D01*
X0011067Y-0026459D02*
Y-0027342D01*
X0011032Y-0026448D02*
Y-0027331D01*
X0010998Y-0026437D02*
Y-0027320D01*
X0010963Y-0026427D02*
Y-0027310D01*
X0010928Y-0026408D02*
Y-0027299D01*
X0010894Y-0026387D02*
Y-0027288D01*
X0010859Y-0026365D02*
Y-0027277D01*
X0010824Y-0026344D02*
Y-0027267D01*
X0010789Y-0026323D02*
Y-0027256D01*
X0010755Y-0026302D02*
Y-0027245D01*
X0010720Y-0026280D02*
Y-0027234D01*
X0010685Y-0026259D02*
Y-0027223D01*
X0010651Y-0026238D02*
Y-0027213D01*
X0010616Y-0026210D02*
Y-0027202D01*
X0010581Y-0026175D02*
Y-0027191D01*
X0010546Y-0026140D02*
Y-0027179D01*
X0010512Y-0026105D02*
Y-0027158D01*
X0010477Y-0026070D02*
Y-0027138D01*
X0010443Y-0026035D02*
Y-0027118D01*
X0010408Y-0026000D02*
Y-0027097D01*
X0010373Y-0025965D02*
Y-0027077D01*
X0010339Y-0025914D02*
Y-0027057D01*
X0010304Y-0025859D02*
Y-0027036D01*
X0010269Y-0025803D02*
Y-0027016D01*
X0010234Y-0025748D02*
Y-0026996D01*
X0010200Y-0025693D02*
Y-0026975D01*
X0010165Y-0025637D02*
Y-0026955D01*
X0010130Y-0025546D02*
Y-0026935D01*
X0010096Y-0025451D02*
Y-0026914D01*
X0010061Y-0025355D02*
Y-0026889D01*
X0010026Y-0025259D02*
Y-0026856D01*
X0009991Y-0025138D02*
Y-0026823D01*
X0009957Y-0025072D02*
Y-0026790D01*
X0009922Y-0025082D02*
Y-0026757D01*
X0009887Y-0025092D02*
Y-0026723D01*
X0009853Y-0025101D02*
Y-0026690D01*
X0009818Y-0025111D02*
Y-0026657D01*
X0009783Y-0025121D02*
Y-0026624D01*
X0009749Y-0025131D02*
Y-0026591D01*
X0009714Y-0025140D02*
Y-0026558D01*
X0009679Y-0025150D02*
Y-0026525D01*
X0009644Y-0025160D02*
Y-0026475D01*
X0009610Y-0025169D02*
Y-0026422D01*
X0009575Y-0025179D02*
Y-0026369D01*
X0009541Y-0025189D02*
Y-0026316D01*
X0009506Y-0025198D02*
Y-0026263D01*
X0009471Y-0025208D02*
Y-0026211D01*
X0009436Y-0025218D02*
Y-0026157D01*
X0009402Y-0025228D02*
Y-0026105D01*
X0009367Y-0025237D02*
Y-0026052D01*
X0009332Y-0025247D02*
Y-0025964D01*
X0009298Y-0025257D02*
Y-0025874D01*
X0009263Y-0025267D02*
Y-0025783D01*
X0009228Y-0025276D02*
Y-0025693D01*
X0009194Y-0025286D02*
Y-0025602D01*
X0009159Y-0025296D02*
Y-0025512D01*
X0012004Y-0019052D02*
X0011732D01*
X0012239Y-0019087D02*
X0011336D01*
X0012414Y-0019121D02*
X0011197D01*
X0012517Y-0019156D02*
X0011058D01*
X0012620Y-0019191D02*
X0010919D01*
X0012724Y-0019225D02*
X0010836D01*
X0012798Y-0019260D02*
X0010768D01*
X0012862Y-0019295D02*
X0010700D01*
X0012925Y-0019330D02*
X0010633D01*
X0012989Y-0019364D02*
X0010565D01*
X0013052Y-0019399D02*
X0010497D01*
X0013113Y-0019433D02*
X0010430D01*
X0013155Y-0019468D02*
X0010380D01*
X0013198Y-0019503D02*
X0010341D01*
X0013240Y-0019537D02*
X0010301D01*
X0013283Y-0019572D02*
X0010261D01*
X0013326Y-0019607D02*
X0010222D01*
X0013368Y-0019642D02*
X0010182D01*
X0013411Y-0019676D02*
X0010143D01*
X0013444Y-0019711D02*
X0010103D01*
X0013474Y-0019746D02*
X0010063D01*
X0013504Y-0019780D02*
X0010024D01*
X0013535Y-0019815D02*
X0009994D01*
X0013565Y-0019850D02*
X0009971D01*
X0011717Y-0019885D02*
X0009948D01*
X0011433Y-0019919D02*
X0009925D01*
X0011323Y-0019954D02*
X0009902D01*
X0011213Y-0019989D02*
X0009880D01*
X0011137Y-0020023D02*
X0009857D01*
X0011079Y-0020058D02*
X0009834D01*
X0011021Y-0020093D02*
X0009811D01*
X0010963Y-0020128D02*
X0009789D01*
X0010905Y-0020162D02*
X0009766D01*
X0010868Y-0020197D02*
X0009743D01*
X0010833Y-0020231D02*
X0009720D01*
X0010799Y-0020266D02*
X0009707D01*
X0010764Y-0020301D02*
X0009696D01*
X0010730Y-0020335D02*
X0009685D01*
X0010695Y-0020370D02*
X0009675D01*
X0010666Y-0020405D02*
X0009664D01*
X0010646Y-0020440D02*
X0009654D01*
X0010626Y-0020474D02*
X0009643D01*
X0010606Y-0020509D02*
X0009632D01*
X0010587Y-0020544D02*
X0009621D01*
X0010567Y-0020578D02*
X0009611D01*
X0010547Y-0020613D02*
X0009600D01*
X0010527Y-0020648D02*
X0009589D01*
X0010511Y-0020683D02*
X0009578D01*
X0010502Y-0020717D02*
X0009568D01*
X0010494Y-0020752D02*
X0009557D01*
X0010485Y-0020787D02*
X0009552D01*
X0010477Y-0020821D02*
X0009551D01*
X0010469Y-0020856D02*
X0009550D01*
X0010460Y-0020891D02*
X0009550D01*
X0010452Y-0020925D02*
X0009548D01*
X0010444Y-0020960D02*
X0009548D01*
X0010435Y-0020995D02*
X0009547D01*
X0010436Y-0021030D02*
X0009546D01*
X0010437Y-0021064D02*
X0009545D01*
X0010439Y-0021099D02*
X0009544D01*
X0010441Y-0021133D02*
X0009543D01*
X0010442Y-0021168D02*
X0009543D01*
X0010444Y-0021203D02*
X0009542D01*
X0010445Y-0021238D02*
X0009541D01*
X0010447Y-0021272D02*
X0009540D01*
X0010448Y-0021307D02*
X0009539D01*
X0010454Y-0021342D02*
X0009541D01*
X0010468Y-0021376D02*
X0009549D01*
X0010482Y-0021411D02*
X0009557D01*
X0010496Y-0021446D02*
X0009565D01*
X0010510Y-0021480D02*
X0009574D01*
X0010524Y-0021515D02*
X0009582D01*
X0010537Y-0021550D02*
X0009590D01*
X0010551Y-0021585D02*
X0009598D01*
X0010570Y-0021619D02*
X0009607D01*
X0010599Y-0021654D02*
X0009615D01*
X0010627Y-0021689D02*
X0009623D01*
X0010656Y-0021723D02*
X0009631D01*
X0010684Y-0021758D02*
X0009640D01*
X0010712Y-0021793D02*
X0009648D01*
X0010741Y-0021828D02*
X0009664D01*
X0010780Y-0021862D02*
X0009683D01*
X0010824Y-0021897D02*
X0009703D01*
X0010867Y-0021931D02*
X0009722D01*
X0010911Y-0021966D02*
X0009741D01*
X0010954Y-0022001D02*
X0009760D01*
X0011001Y-0022035D02*
X0009780D01*
X0011059Y-0022070D02*
X0009799D01*
X0011119Y-0022105D02*
X0009818D01*
X0011178Y-0022140D02*
X0009837D01*
X0011237Y-0022174D02*
X0009856D01*
X0011303Y-0022209D02*
X0009883D01*
X0011374Y-0022244D02*
X0009916D01*
X0011445Y-0022278D02*
X0009948D01*
X0011516Y-0022313D02*
X0009981D01*
X0011591Y-0022348D02*
X0010013D01*
X0011668Y-0022383D02*
X0010046D01*
X0011746Y-0022417D02*
X0010078D01*
X0011826Y-0022452D02*
X0010111D01*
X0011905Y-0022487D02*
X0010143D01*
X0011983Y-0022521D02*
X0010181D01*
X0012061Y-0022556D02*
X0010229D01*
X0012139Y-0022591D02*
X0010277D01*
X0012217Y-0022626D02*
X0010325D01*
X0012295Y-0022660D02*
X0010372D01*
X0012372Y-0022695D02*
X0010420D01*
X0012443Y-0022730D02*
X0010468D01*
X0012514Y-0022764D02*
X0010516D01*
X0012585Y-0022799D02*
X0010574D01*
X0012656Y-0022833D02*
X0010636D01*
X0012727Y-0022868D02*
X0010699D01*
X0012798Y-0022903D02*
X0010761D01*
X0012863Y-0022938D02*
X0010824D01*
X0012920Y-0022972D02*
X0010886D01*
X0012976Y-0023007D02*
X0010949D01*
X0013033Y-0023042D02*
X0011022D01*
X0013089Y-0023076D02*
X0011095D01*
X0013146Y-0023111D02*
X0011169D01*
X0013202Y-0023146D02*
X0011241D01*
X0013259Y-0023181D02*
X0011318D01*
X0013304Y-0023215D02*
X0011398D01*
X0013344Y-0023250D02*
X0011478D01*
X0013384Y-0023285D02*
X0011559D01*
X0013424Y-0023319D02*
X0011637D01*
X0013464Y-0023354D02*
X0011716D01*
X0013504Y-0023389D02*
X0011797D01*
X0013544Y-0023423D02*
X0011871D01*
X0013585Y-0023458D02*
X0011945D01*
X0013625Y-0023493D02*
X0012019D01*
X0013658Y-0023528D02*
X0012093D01*
X0013683Y-0023562D02*
X0012166D01*
X0013709Y-0023597D02*
X0012231D01*
X0013734Y-0023631D02*
X0012296D01*
X0013760Y-0023666D02*
X0012361D01*
X0013785Y-0023701D02*
X0012426D01*
X0013811Y-0023736D02*
X0012491D01*
X0013837Y-0023770D02*
X0012542D01*
X0013862Y-0023805D02*
X0012590D01*
X0013888Y-0023840D02*
X0012639D01*
X0013913Y-0023874D02*
X0012687D01*
X0013935Y-0023909D02*
X0012736D01*
X0013948Y-0023944D02*
X0012785D01*
X0013961Y-0023978D02*
X0012821D01*
X0013974Y-0024013D02*
X0012853D01*
X0013987Y-0024048D02*
X0012885D01*
X0014001Y-0024083D02*
X0012917D01*
X0014014Y-0024117D02*
X0012950D01*
X0014027Y-0024152D02*
X0012982D01*
X0014041Y-0024187D02*
X0013014D01*
X0014054Y-0024221D02*
X0013042D01*
X0014067Y-0024256D02*
X0013059D01*
X0014080Y-0024291D02*
X0013077D01*
X0014094Y-0024326D02*
X0013095D01*
X0014107Y-0024360D02*
X0013113D01*
X0014113Y-0024395D02*
X0013130D01*
X0014116Y-0024430D02*
X0013148D01*
X0014120Y-0024464D02*
X0013166D01*
X0014123Y-0024499D02*
X0013183D01*
X0014127Y-0024533D02*
X0013200D01*
X0014130Y-0024569D02*
X0013206D01*
X0014134Y-0024603D02*
X0013212D01*
X0014137Y-0024638D02*
X0013218D01*
X0014141Y-0024672D02*
X0013224D01*
X0014144Y-0024707D02*
X0013230D01*
X0014148Y-0024742D02*
X0013235D01*
X0014151Y-0024776D02*
X0013241D01*
X0014155Y-0024811D02*
X0013247D01*
X0014158Y-0024846D02*
X0013253D01*
X0014162Y-0024881D02*
X0013259D01*
X0014165Y-0024915D02*
X0013265D01*
X0014168Y-0024950D02*
X0013266D01*
X0014163Y-0024985D02*
X0013262D01*
X0014157Y-0025019D02*
X0013258D01*
X0014152Y-0025054D02*
X0013255D01*
X0009977Y-0025089D02*
X0009898D01*
X0009987Y-0025124D02*
X0009774D01*
X0009997Y-0025158D02*
X0009650D01*
X0010007Y-0025193D02*
X0009526D01*
X0010017Y-0025228D02*
X0009403D01*
X0010027Y-0025262D02*
X0009280D01*
X0010040Y-0025297D02*
X0009155D01*
X0010052Y-0025331D02*
X0009141D01*
X0010065Y-0025366D02*
X0009143D01*
X0010078Y-0025401D02*
X0009146D01*
X0010090Y-0025436D02*
X0009149D01*
X0010103Y-0025470D02*
X0009151D01*
X0010115Y-0025505D02*
X0009156D01*
X0010128Y-0025540D02*
X0009170D01*
X0010141Y-0025574D02*
X0009183D01*
X0010153Y-0025609D02*
X0009196D01*
X0010169Y-0025644D02*
X0009209D01*
X0010191Y-0025679D02*
X0009223D01*
X0010213Y-0025713D02*
X0009236D01*
X0010234Y-0025748D02*
X0009249D01*
X0010256Y-0025783D02*
X0009263D01*
X0010278Y-0025817D02*
X0009276D01*
X0010300Y-0025852D02*
X0009289D01*
X0010321Y-0025887D02*
X0009303D01*
X0010343Y-0025921D02*
X0009316D01*
X0010365Y-0025956D02*
X0009329D01*
X0010399Y-0025991D02*
X0009343D01*
X0010433Y-0026026D02*
X0009356D01*
X0010468Y-0026060D02*
X0009372D01*
X0010502Y-0026095D02*
X0009395D01*
X0010536Y-0026130D02*
X0009418D01*
X0010570Y-0026164D02*
X0009441D01*
X0010605Y-0026199D02*
X0009463D01*
X0010644Y-0026234D02*
X0009486D01*
X0010701Y-0026269D02*
X0009509D01*
X0010757Y-0026303D02*
X0009532D01*
X0010814Y-0026338D02*
X0009555D01*
X0010870Y-0026372D02*
X0009577D01*
X0010927Y-0026407D02*
X0009600D01*
X0011012Y-0026442D02*
X0009623D01*
X0011124Y-0026476D02*
X0009646D01*
X0011236Y-0026511D02*
X0009669D01*
X0011462Y-0026546D02*
X0009702D01*
X0013507Y-0026581D02*
X0009738D01*
X0013480Y-0026615D02*
X0009774D01*
X0013453Y-0026650D02*
X0009811D01*
X0013418Y-0026685D02*
X0009847D01*
X0013373Y-0026719D02*
X0009883D01*
X0013328Y-0026754D02*
X0009920D01*
X0013282Y-0026789D02*
X0009956D01*
X0013237Y-0026824D02*
X0009992D01*
X0013191Y-0026858D02*
X0010029D01*
X0013146Y-0026893D02*
X0010065D01*
X0013101Y-0026928D02*
X0010119D01*
X0013056Y-0026962D02*
X0010178D01*
X0013010Y-0026997D02*
X0010237D01*
X0012965Y-0027031D02*
X0010296D01*
X0012900Y-0027067D02*
X0010355D01*
X0012819Y-0027101D02*
X0010414D01*
X0012738Y-0027136D02*
X0010473D01*
X0012657Y-0027170D02*
X0010533D01*
X0012577Y-0027205D02*
X0010627D01*
X0012496Y-0027240D02*
X0010739D01*
X0012415Y-0027274D02*
X0010850D01*
X0012287Y-0027309D02*
X0010961D01*
X0012065Y-0027344D02*
X0011073D01*
X0013843Y-0020237D02*
Y-0020317D01*
X0013808Y-0020181D02*
Y-0020339D01*
X0013773Y-0020126D02*
Y-0020361D01*
X0013739Y-0020070D02*
Y-0020383D01*
X0013704Y-0020014D02*
Y-0020405D01*
X0013669Y-0019969D02*
Y-0020427D01*
X0013635Y-0019930D02*
Y-0020450D01*
X0013600Y-0019890D02*
Y-0020472D01*
X0013565Y-0019850D02*
Y-0020495D01*
X0013530Y-0019810D02*
Y-0020517D01*
X0013496Y-0019770D02*
Y-0020540D01*
X0013461Y-0019731D02*
Y-0020562D01*
X0013426Y-0019691D02*
Y-0020584D01*
X0013392Y-0019661D02*
Y-0020606D01*
X0013357Y-0019633D02*
Y-0020628D01*
X0013322Y-0019604D02*
Y-0020651D01*
X0013287Y-0019576D02*
Y-0020673D01*
X0008922Y-0022662D02*
X0008077D01*
X0008924Y-0022696D02*
X0008082D01*
X0008926Y-0022731D02*
X0008087D01*
X0008929Y-0022766D02*
X0008091D01*
X0008931Y-0022800D02*
X0008095D01*
X0008933Y-0022835D02*
X0008100D01*
X0008936Y-0022870D02*
X0008104D01*
X0008939Y-0022905D02*
X0008108D01*
X0008941Y-0022939D02*
X0008110D01*
X0008943Y-0022974D02*
X0008112D01*
X0008946Y-0023009D02*
X0008114D01*
X0008948Y-0023043D02*
X0008116D01*
X0008950Y-0023078D02*
X0008119D01*
X0008953Y-0023113D02*
X0008120D01*
X0008956Y-0023148D02*
X0008120D01*
X0008958Y-0023182D02*
X0008120D01*
X0008960Y-0023217D02*
X0008120D01*
X0008963Y-0023252D02*
X0008120D01*
X0008965Y-0023286D02*
X0008120D01*
X0008968Y-0023321D02*
X0008120D01*
X0008970Y-0023356D02*
X0008119D01*
X0008972Y-0023390D02*
X0008116D01*
X0008969Y-0023425D02*
X0008114D01*
X0008963Y-0023460D02*
X0008112D01*
X0008958Y-0023494D02*
X0008109D01*
X0008952Y-0023529D02*
X0008107D01*
X0008946Y-0023564D02*
X0008104D01*
X0008941Y-0023598D02*
X0008100D01*
X0008935Y-0023633D02*
X0008095D01*
X0008930Y-0023668D02*
X0008091D01*
X0008924Y-0023703D02*
X0008086D01*
X0008919Y-0023737D02*
X0008081D01*
X0008913Y-0023772D02*
X0008076D01*
X0008907Y-0023807D02*
X0008070D01*
X0008902Y-0023841D02*
X0008063D01*
X0008896Y-0023876D02*
X0008056D01*
X0008891Y-0023911D02*
X0008049D01*
X0008885Y-0023945D02*
X0008042D01*
X0008880Y-0023980D02*
X0008035D01*
X0008874Y-0024015D02*
X0008025D01*
X0008869Y-0024050D02*
X0008016D01*
X0008863Y-0024084D02*
X0008007D01*
X0008857Y-0024119D02*
X0007998D01*
X0008852Y-0024154D02*
X0007989D01*
X0008846Y-0024188D02*
X0007979D01*
X0008841Y-0024223D02*
X0007967D01*
X0008835Y-0024258D02*
X0007956D01*
X0008830Y-0024293D02*
X0007944D01*
X0008824Y-0024327D02*
X0007932D01*
X0008819Y-0024362D02*
X0007920D01*
X0008813Y-0024396D02*
X0007907D01*
X0008807Y-0024431D02*
X0007894D01*
X0008802Y-0024466D02*
X0007880D01*
X0008792Y-0024500D02*
X0007865D01*
X0008775Y-0024535D02*
X0007852D01*
X0008758Y-0024570D02*
X0007837D01*
X0008741Y-0024605D02*
X0007821D01*
X0008724Y-0024639D02*
X0007804D01*
X0008707Y-0024674D02*
X0007787D01*
X0008689Y-0024709D02*
X0007771D01*
X0008672Y-0024743D02*
X0007754D01*
X0008655Y-0024778D02*
X0007736D01*
X0008638Y-0024813D02*
X0007717D01*
X0008621Y-0024848D02*
X0007697D01*
X0008604Y-0024882D02*
X0007678D01*
X0008587Y-0024917D02*
X0007658D01*
X0008570Y-0024952D02*
X0007638D01*
X0008553Y-0024986D02*
X0007616D01*
X0008535Y-0025021D02*
X0007594D01*
X0008519Y-0025056D02*
X0007572D01*
X0008501Y-0025091D02*
X0007549D01*
X0008484Y-0025125D02*
X0007526D01*
X0008467Y-0025160D02*
X0007501D01*
X0008450Y-0025194D02*
X0007475D01*
X0008433Y-0025229D02*
X0007450D01*
X0008416Y-0025264D02*
X0007424D01*
X0008399Y-0025298D02*
X0007397D01*
X0008381Y-0025333D02*
X0007369D01*
X0008365Y-0025368D02*
X0007340D01*
X0008347Y-0025403D02*
X0007311D01*
X0008330Y-0025437D02*
X0007283D01*
X0008303Y-0025472D02*
X0007251D01*
X0008274Y-0025507D02*
X0007218D01*
X0008245Y-0025541D02*
X0007185D01*
X0008215Y-0025576D02*
X0007153D01*
X0008186Y-0025611D02*
X0007119D01*
X0008157Y-0025646D02*
X0007081D01*
X0008128Y-0025680D02*
X0007044D01*
X0008099Y-0025715D02*
X0007007D01*
X0008070Y-0025750D02*
X0006968D01*
X0008041Y-0025784D02*
X0006926D01*
X0008011Y-0025819D02*
X0006884D01*
X0007982Y-0025854D02*
X0006842D01*
X0007953Y-0025888D02*
X0006797D01*
X0007924Y-0025923D02*
X0006750D01*
X0007894Y-0025958D02*
X0006703D01*
X0007865Y-0025993D02*
X0006656D01*
X0007836Y-0026027D02*
X0006601D01*
X0007807Y-0026062D02*
X0006546D01*
X0007778Y-0026096D02*
X0006492D01*
X0007749Y-0026131D02*
X0006431D01*
X0007720Y-0026166D02*
X0006368D01*
X0007691Y-0026201D02*
X0006306D01*
X0007648Y-0026235D02*
X0006233D01*
X0007602Y-0026270D02*
X0006161D01*
X0007555Y-0026305D02*
X0006083D01*
X0007508Y-0026339D02*
X0005997D01*
X0007461Y-0026374D02*
X0005908D01*
X0007414Y-0026409D02*
X0005803D01*
X0007367Y-0026443D02*
X0005691D01*
X0007320Y-0026478D02*
X0005553D01*
X0007274Y-0026513D02*
X0005380D01*
X0007227Y-0026548D02*
X0005129D01*
X0007180Y-0026582D02*
X0004669D01*
X0007133Y-0026617D02*
X0004670D01*
X0007087Y-0026652D02*
X0004670D01*
X0007040Y-0026686D02*
X0004671D01*
X0006993Y-0026721D02*
X0004672D01*
X0006946Y-0026756D02*
X0004672D01*
X0006898Y-0026791D02*
X0004673D01*
X0006827Y-0026825D02*
X0004674D01*
X0006756Y-0026860D02*
X0004674D01*
X0006685Y-0026894D02*
X0004675D01*
X0006615Y-0026929D02*
X0004675D01*
X0006544Y-0026964D02*
X0004676D01*
X0006473Y-0026998D02*
X0004676D01*
X0006402Y-0027033D02*
X0004677D01*
X0006331Y-0027068D02*
X0004678D01*
X0006261Y-0027103D02*
X0004678D01*
X0006190Y-0027137D02*
X0004679D01*
X0006066Y-0027172D02*
X0004679D01*
X0005908Y-0027207D02*
X0004680D01*
X0005750Y-0027241D02*
X0004680D01*
X0005592Y-0027276D02*
X0004681D01*
X0005433Y-0027311D02*
X0004681D01*
X0004969Y-0027346D02*
X0004682D01*
X0004645D02*
X0004510D01*
X0001505Y-0022999D02*
X0001498Y-0023220D01*
X0001525Y-0022782D02*
X0001505Y-0022999D01*
X0001560Y-0022570D02*
X0001525Y-0022782D01*
X0001608Y-0022361D02*
X0001560Y-0022570D01*
X0001668Y-0022158D02*
X0001608Y-0022361D01*
X0001739Y-0021960D02*
X0001668Y-0022158D01*
X0001824Y-0021769D02*
X0001739Y-0021960D01*
X0001919Y-0021583D02*
X0001824Y-0021769D01*
X0002025Y-0021405D02*
X0001919Y-0021583D01*
X0002142Y-0021234D02*
X0002025Y-0021405D01*
X0002269Y-0021071D02*
X0002142Y-0021234D01*
X0002406Y-0020916D02*
X0002269Y-0021071D01*
X0002550Y-0020770D02*
X0002406Y-0020916D01*
X0002706Y-0020633D02*
X0002550Y-0020770D01*
X0002868Y-0020506D02*
X0002706Y-0020633D01*
X0003039Y-0020389D02*
X0002868Y-0020506D01*
X0003217Y-0020283D02*
X0003039Y-0020389D01*
X0003403Y-0020188D02*
X0003217Y-0020283D01*
X0003595Y-0020106D02*
X0003403Y-0020188D01*
X0003794Y-0020034D02*
X0003595Y-0020106D01*
X0003998Y-0019976D02*
X0003794Y-0020034D01*
X0004209Y-0019929D02*
X0003998Y-0019976D01*
X0004424Y-0019898D02*
X0004209Y-0019929D01*
X0004643Y-0019878D02*
X0004424Y-0019898D01*
X0004866Y-0019876D02*
X0004643Y-0019878D01*
X0004866Y-0019876D02*
X0005088Y-0019887D01*
X0005306Y-0019913D01*
X0005517Y-0019951D01*
X0005726Y-0020003D01*
X0005927Y-0020068D01*
X0006122Y-0020145D01*
X0006311Y-0020235D01*
X0006494Y-0020335D01*
X0006668Y-0020446D01*
X0006835Y-0020569D01*
X0006994Y-0020700D01*
X0007144Y-0020842D01*
X0007285Y-0020992D01*
X0007417Y-0021151D01*
X0007538Y-0021318D01*
X0007650Y-0021493D01*
X0007750Y-0021675D01*
X0007840Y-0021864D01*
X0007919Y-0022058D01*
X0007985Y-0022259D01*
X0008038Y-0022465D01*
X0008080Y-0022675D01*
X0008107Y-0022891D01*
X0008120Y-0023109D01*
Y-0023330D01*
X0008106Y-0023547D01*
X0008079Y-0023761D01*
X0008037Y-0023972D01*
X0007983Y-0024177D01*
X0007916Y-0024377D01*
X0007837Y-0024572D01*
X0007746Y-0024760D01*
X0007645Y-0024942D01*
X0007532Y-0025117D01*
X0007410Y-0025283D01*
X0007278Y-0025443D01*
X0007136Y-0025594D01*
X0006985Y-0025735D01*
X0006825Y-0025868D01*
X0006659Y-0025991D01*
X0006483Y-0026102D01*
X0006302Y-0026203D01*
X0006113Y-0026293D01*
X0005919Y-0026371D01*
X0005717Y-0026437D01*
X0005511Y-0026489D01*
X0005301Y-0026528D01*
X0005087Y-0026553D01*
X0004866Y-0026565D01*
X0004669Y-0026560D02*
X0004866Y-0026565D01*
X0004669Y-0026560D02*
X0004683Y-0027366D01*
X0005423Y-0027313D02*
X0004683Y-0027366D01*
X0006162Y-0027151D02*
X0005423Y-0027313D01*
X0006902Y-0026789D02*
X0006162Y-0027151D01*
X0007683Y-0026210D02*
X0006902Y-0026789D01*
X0008328Y-0025443D02*
X0007683Y-0026210D01*
X0008798Y-0024488D02*
X0008328Y-0025443D01*
X0008973Y-0023399D02*
X0008798Y-0024488D01*
X0008906Y-0022431D02*
X0008973Y-0023399D01*
X0008650Y-0021610D02*
X0008906Y-0022431D01*
X0008112Y-0020696D02*
X0008650Y-0021610D01*
X0007372Y-0019983D02*
X0008112Y-0020696D01*
X0006633Y-0019486D02*
X0007372Y-0019983D01*
X0005746Y-0019176D02*
X0006633Y-0019486D01*
X0004724Y-0019082D02*
X0005746Y-0019176D01*
X0004724Y-0019082D02*
X0003809Y-0019217D01*
X0002854Y-0019580D01*
X0001993Y-0020186D01*
X0001402Y-0020871D01*
X0000971Y-0021665D01*
X0000689Y-0022592D01*
X0000648Y-0023561D01*
X0000864Y-0024543D01*
X0001348Y-0025551D01*
X0002141Y-0026385D01*
X0002934Y-0026923D01*
X0003849Y-0027246D01*
X0004645Y-0027366D01*
Y-0026561D02*
Y-0027366D01*
X0004427Y-0026542D02*
X0004645Y-0026561D01*
X0004214Y-0026509D02*
X0004427Y-0026542D01*
X0004006Y-0026464D02*
X0004214Y-0026509D01*
X0003802Y-0026405D02*
X0004006Y-0026464D01*
X0003604Y-0026333D02*
X0003802Y-0026405D01*
X0003413Y-0026250D02*
X0003604Y-0026333D01*
X0003227Y-0026154D02*
X0003413Y-0026250D01*
X0003049Y-0026048D02*
X0003227Y-0026154D01*
X0002877Y-0025931D02*
X0003049Y-0026048D01*
X0002714Y-0025803D02*
X0002877Y-0025931D01*
X0002558Y-0025666D02*
X0002714Y-0025803D01*
X0002413Y-0025520D02*
X0002558Y-0025666D01*
X0002276Y-0025365D02*
X0002413Y-0025520D01*
X0002149Y-0025202D02*
X0002276Y-0025365D01*
X0002031Y-0025030D02*
X0002149Y-0025202D01*
X0001924Y-0024852D02*
X0002031Y-0025030D01*
X0001828Y-0024667D02*
X0001924Y-0024852D01*
X0001743Y-0024475D02*
X0001828Y-0024667D01*
X0001670Y-0024278D02*
X0001743Y-0024475D01*
X0001609Y-0024075D02*
X0001670Y-0024278D01*
X0001561Y-0023867D02*
X0001609Y-0024075D01*
X0001526Y-0023655D02*
X0001561Y-0023867D01*
X0001506Y-0023439D02*
X0001526Y-0023655D01*
X0001498Y-0023220D02*
X0001506Y-0023439D01*
X0008960Y-0023217D02*
Y-0023478D01*
X0008926Y-0022721D02*
Y-0023694D01*
X0008891Y-0022384D02*
Y-0023910D01*
X0008856Y-0022273D02*
Y-0024126D01*
X0008822Y-0022161D02*
Y-0024343D01*
X0008787Y-0022050D02*
Y-0024511D01*
X0008752Y-0021938D02*
Y-0024581D01*
X0008717Y-0021826D02*
Y-0024652D01*
X0008683Y-0021715D02*
Y-0024722D01*
X0008648Y-0021606D02*
Y-0024793D01*
X0008613Y-0021548D02*
Y-0024863D01*
X0008579Y-0021489D02*
Y-0024933D01*
X0008544Y-0021430D02*
Y-0025004D01*
X0008509Y-0021371D02*
Y-0025074D01*
X0008475Y-0021312D02*
Y-0025144D01*
X0008440Y-0021253D02*
Y-0025215D01*
X0008405Y-0021194D02*
Y-0025285D01*
X0008370Y-0021135D02*
Y-0025356D01*
X0008336Y-0021076D02*
Y-0025426D01*
X0008301Y-0021018D02*
Y-0025474D01*
X0008267Y-0020959D02*
Y-0025516D01*
X0008232Y-0020900D02*
Y-0025557D01*
X0008197Y-0020841D02*
Y-0025598D01*
X0008162Y-0020782D02*
Y-0025639D01*
X0008128Y-0020723D02*
Y-0025681D01*
X0008093Y-0023649D02*
Y-0025722D01*
X0008058Y-0023863D02*
Y-0025763D01*
X0008024Y-0024022D02*
Y-0025804D01*
X0007989Y-0024153D02*
Y-0025846D01*
X0007954Y-0024261D02*
Y-0025887D01*
X0007920Y-0024365D02*
Y-0025928D01*
X0007885Y-0024453D02*
Y-0025969D01*
X0007850Y-0024539D02*
Y-0026011D01*
X0007815Y-0024616D02*
Y-0026052D01*
X0007781Y-0024688D02*
Y-0026093D01*
X0007746Y-0024760D02*
Y-0026135D01*
X0007711Y-0024822D02*
Y-0026176D01*
X0007677Y-0024884D02*
Y-0026215D01*
X0007642Y-0024946D02*
Y-0026240D01*
X0007607Y-0025000D02*
Y-0026266D01*
X0007572Y-0025054D02*
Y-0026291D01*
X0007538Y-0025108D02*
Y-0026317D01*
X0007503Y-0025157D02*
Y-0026343D01*
X0007469Y-0025204D02*
Y-0026369D01*
X0007434Y-0025251D02*
Y-0026394D01*
X0007399Y-0025296D02*
Y-0026420D01*
X0007365Y-0025339D02*
Y-0026446D01*
X0007330Y-0025380D02*
Y-0026471D01*
X0007295Y-0025422D02*
Y-0026497D01*
X0007260Y-0025462D02*
Y-0026523D01*
X0007226Y-0025499D02*
Y-0026548D01*
X0007191Y-0025536D02*
Y-0026574D01*
X0007156Y-0025573D02*
Y-0026600D01*
X0007122Y-0025608D02*
Y-0026626D01*
X0007087Y-0025640D02*
Y-0026652D01*
X0007052Y-0025672D02*
Y-0026677D01*
X0007017Y-0025705D02*
Y-0026703D01*
X0006983Y-0025737D02*
Y-0026728D01*
X0006948Y-0025766D02*
Y-0026754D01*
X0006913Y-0025794D02*
Y-0026780D01*
X0006879Y-0025823D02*
Y-0026800D01*
X0006844Y-0025852D02*
Y-0026817D01*
X0006809Y-0025879D02*
Y-0026834D01*
X0006774Y-0025905D02*
Y-0026851D01*
X0006740Y-0025930D02*
Y-0026868D01*
X0006705Y-0025956D02*
Y-0026885D01*
X0006670Y-0025982D02*
Y-0026902D01*
X0006636Y-0026005D02*
Y-0026919D01*
X0006601Y-0026027D02*
Y-0026936D01*
X0006567Y-0026049D02*
Y-0026953D01*
X0006532Y-0026071D02*
Y-0026970D01*
X0006497Y-0026093D02*
Y-0026987D01*
X0006462Y-0026114D02*
Y-0027004D01*
X0006428Y-0026133D02*
Y-0027021D01*
X0006393Y-0026152D02*
Y-0027038D01*
X0006358Y-0026172D02*
Y-0027055D01*
X0006324Y-0026191D02*
Y-0027072D01*
X0006289Y-0026209D02*
Y-0027089D01*
X0006254Y-0026226D02*
Y-0027106D01*
X0006219Y-0026242D02*
Y-0027123D01*
X0006185Y-0026259D02*
Y-0027140D01*
X0006150Y-0026275D02*
Y-0027154D01*
X0006115Y-0026292D02*
Y-0027161D01*
X0006081Y-0026306D02*
Y-0027169D01*
X0006046Y-0026320D02*
Y-0027176D01*
X0006011Y-0026333D02*
Y-0027184D01*
X0005977Y-0026348D02*
Y-0027192D01*
X0005942Y-0026361D02*
Y-0027199D01*
X0005907Y-0026374D02*
Y-0027207D01*
X0005872Y-0026386D02*
Y-0027215D01*
X0005838Y-0026397D02*
Y-0027222D01*
X0005803Y-0026409D02*
Y-0027230D01*
X0005769Y-0026420D02*
Y-0027237D01*
X0005734Y-0026431D02*
Y-0027245D01*
X0005699Y-0026441D02*
Y-0027252D01*
X0005664Y-0026450D02*
Y-0027260D01*
X0005630Y-0026459D02*
Y-0027268D01*
X0005595Y-0026468D02*
Y-0027275D01*
X0005560Y-0026476D02*
Y-0027283D01*
X0005526Y-0026485D02*
Y-0027291D01*
X0005491Y-0026493D02*
Y-0027298D01*
X0005456Y-0026499D02*
Y-0027306D01*
X0005422Y-0026505D02*
Y-0027313D01*
X0005387Y-0026511D02*
Y-0027316D01*
X0005352Y-0026518D02*
Y-0027318D01*
X0005317Y-0026524D02*
Y-0027321D01*
X0005283Y-0026530D02*
Y-0027323D01*
X0005248Y-0026533D02*
Y-0027326D01*
X0005213Y-0026538D02*
Y-0027328D01*
X0005179Y-0026542D02*
Y-0027331D01*
X0005144Y-0026546D02*
Y-0027333D01*
X0005109Y-0026550D02*
Y-0027335D01*
X0005074Y-0026553D02*
Y-0027338D01*
X0005040Y-0026555D02*
Y-0027341D01*
X0005005Y-0026557D02*
Y-0027343D01*
X0004970Y-0026559D02*
Y-0027345D01*
X0004936Y-0026561D02*
Y-0027348D01*
X0004901Y-0026563D02*
Y-0027350D01*
X0004867Y-0026564D02*
Y-0027353D01*
X0004831Y-0026563D02*
Y-0027355D01*
X0004797Y-0026563D02*
Y-0027358D01*
X0004762Y-0026562D02*
Y-0027360D01*
X0004728Y-0026561D02*
Y-0027363D01*
X0004693Y-0026560D02*
Y-0027365D01*
X0004658Y-0019091D02*
Y-0019878D01*
X0004624Y-0026559D02*
Y-0027363D01*
X0004589Y-0026556D02*
Y-0027357D01*
X0004554Y-0026553D02*
Y-0027352D01*
X0004519Y-0026550D02*
Y-0027347D01*
X0004485Y-0026546D02*
Y-0027342D01*
X0004450Y-0026544D02*
Y-0027337D01*
X0004415Y-0026540D02*
Y-0027331D01*
X0004381Y-0026535D02*
Y-0027326D01*
X0004346Y-0026529D02*
Y-0027321D01*
X0004311Y-0026524D02*
Y-0027315D01*
X0004276Y-0026519D02*
Y-0027310D01*
X0004242Y-0026513D02*
Y-0027305D01*
X0004207Y-0026508D02*
Y-0027300D01*
X0004172Y-0026500D02*
Y-0027294D01*
X0004138Y-0026493D02*
Y-0027289D01*
X0004103Y-0026485D02*
Y-0027284D01*
X0004069Y-0026478D02*
Y-0027279D01*
X0004034Y-0026470D02*
Y-0027274D01*
X0003999Y-0026462D02*
Y-0027268D01*
X0003964Y-0026452D02*
Y-0027263D01*
X0003930Y-0026442D02*
Y-0027258D01*
X0003895Y-0026431D02*
Y-0027252D01*
X0003860Y-0026422D02*
Y-0027247D01*
X0003826Y-0026411D02*
Y-0027237D01*
X0003791Y-0026401D02*
Y-0027225D01*
X0003756Y-0026388D02*
Y-0027213D01*
X0003721Y-0026376D02*
Y-0027200D01*
X0003687Y-0026363D02*
Y-0027188D01*
X0003652Y-0026350D02*
Y-0027176D01*
X0003617Y-0026338D02*
Y-0027164D01*
X0003583Y-0026324D02*
Y-0027152D01*
X0003548Y-0026309D02*
Y-0027139D01*
X0003513Y-0026293D02*
Y-0027127D01*
X0003479Y-0026278D02*
Y-0027115D01*
X0003444Y-0026263D02*
Y-0027103D01*
X0003409Y-0026248D02*
Y-0027091D01*
X0003374Y-0026230D02*
Y-0027078D01*
X0003340Y-0026212D02*
Y-0027066D01*
X0003305Y-0026194D02*
Y-0027054D01*
X0003270Y-0026177D02*
Y-0027041D01*
X0003236Y-0026159D02*
Y-0027029D01*
X0003201Y-0026139D02*
Y-0027017D01*
X0003166Y-0026118D02*
Y-0027005D01*
X0003131Y-0026097D02*
Y-0026993D01*
X0003097Y-0026077D02*
Y-0026980D01*
X0003062Y-0026056D02*
Y-0026968D01*
X0003028Y-0026033D02*
Y-0026956D01*
X0002993Y-0026010D02*
Y-0026944D01*
X0002958Y-0025986D02*
Y-0026931D01*
X0002924Y-0025962D02*
Y-0026916D01*
X0002889Y-0025939D02*
Y-0026892D01*
X0002854Y-0025913D02*
Y-0026869D01*
X0002819Y-0025885D02*
Y-0026845D01*
X0002785Y-0025858D02*
Y-0026822D01*
X0002750Y-0025831D02*
Y-0026798D01*
X0002715Y-0025804D02*
Y-0026774D01*
X0002681Y-0025774D02*
Y-0026751D01*
X0002646Y-0025743D02*
Y-0026728D01*
X0002611Y-0025713D02*
Y-0026704D01*
X0002576Y-0025682D02*
Y-0026680D01*
X0002542Y-0025650D02*
Y-0026657D01*
X0002507Y-0025615D02*
Y-0026633D01*
X0002472Y-0025580D02*
Y-0026610D01*
X0002438Y-0025544D02*
Y-0026586D01*
X0002403Y-0025508D02*
Y-0026563D01*
X0002369Y-0025469D02*
Y-0026539D01*
X0002333Y-0025430D02*
Y-0026516D01*
X0002299Y-0025391D02*
Y-0026492D01*
X0002264Y-0025350D02*
Y-0026469D01*
X0002230Y-0025306D02*
Y-0026445D01*
X0002195Y-0025261D02*
Y-0026422D01*
X0002160Y-0025216D02*
Y-0026398D01*
X0002126Y-0025168D02*
Y-0026369D01*
X0002091Y-0025117D02*
Y-0026332D01*
X0002056Y-0025067D02*
Y-0026296D01*
X0002021Y-0025015D02*
Y-0026259D01*
X0001987Y-0024957D02*
Y-0026223D01*
X0001952Y-0024899D02*
Y-0026186D01*
X0001917Y-0024840D02*
Y-0026150D01*
X0001883Y-0024773D02*
Y-0026113D01*
X0001848Y-0024706D02*
Y-0026077D01*
X0001813Y-0024635D02*
Y-0026041D01*
X0001778Y-0024556D02*
Y-0026004D01*
X0001744Y-0024478D02*
Y-0025967D01*
X0001709Y-0024384D02*
Y-0025931D01*
X0001674Y-0024290D02*
Y-0025894D01*
X0001640Y-0024178D02*
Y-0025858D01*
X0001605Y-0024060D02*
Y-0025821D01*
X0001570Y-0023909D02*
Y-0025785D01*
X0001536Y-0023715D02*
Y-0025748D01*
X0001501Y-0023317D02*
Y-0025712D01*
X0001466Y-0020796D02*
Y-0025676D01*
X0001431Y-0020836D02*
Y-0025639D01*
X0001397Y-0020879D02*
Y-0025602D01*
X0001362Y-0020943D02*
Y-0025566D01*
X0001328Y-0021007D02*
Y-0025509D01*
X0001293Y-0021071D02*
Y-0025436D01*
X0001258Y-0021135D02*
Y-0025364D01*
X0001223Y-0021199D02*
Y-0025292D01*
X0001189Y-0021263D02*
Y-0025219D01*
X0001154Y-0021326D02*
Y-0025147D01*
X0001119Y-0021391D02*
Y-0025075D01*
X0001085Y-0021454D02*
Y-0025003D01*
X0001050Y-0021519D02*
Y-0024930D01*
X0001015Y-0021582D02*
Y-0024858D01*
X0000981Y-0021646D02*
Y-0024786D01*
X0000946Y-0021746D02*
Y-0024714D01*
X0000911Y-0021860D02*
Y-0024641D01*
X0000876Y-0021974D02*
Y-0024569D01*
X0000842Y-0022089D02*
Y-0024443D01*
X0000807Y-0022203D02*
Y-0024285D01*
X0000772Y-0022317D02*
Y-0024127D01*
X0000738Y-0022431D02*
Y-0023969D01*
X0000703Y-0022545D02*
Y-0023811D01*
X0000668Y-0023077D02*
Y-0023654D01*
X0004793Y-0019088D02*
X0004680D01*
X0005169Y-0019123D02*
X0004444D01*
X0005544Y-0019157D02*
X0004208D01*
X0005791Y-0019192D02*
X0003972D01*
X0005891Y-0019227D02*
X0003781D01*
X0005991Y-0019262D02*
X0003689D01*
X0006090Y-0019296D02*
X0003598D01*
X0006189Y-0019331D02*
X0003507D01*
X0006289Y-0019366D02*
X0003415D01*
X0006389Y-0019400D02*
X0003324D01*
X0006488Y-0019435D02*
X0003233D01*
X0006587Y-0019470D02*
X0003142D01*
X0006661Y-0019504D02*
X0003050D01*
X0006713Y-0019539D02*
X0002959D01*
X0006764Y-0019574D02*
X0002868D01*
X0006815Y-0019609D02*
X0002812D01*
X0006867Y-0019643D02*
X0002763D01*
X0006919Y-0019678D02*
X0002713D01*
X0006970Y-0019713D02*
X0002664D01*
X0007022Y-0019747D02*
X0002615D01*
X0007073Y-0019782D02*
X0002566D01*
X0007125Y-0019817D02*
X0002517D01*
X0007176Y-0019852D02*
X0002467D01*
X0004550Y-0019886D02*
X0002418D01*
X0004264Y-0019921D02*
X0002369D01*
X0004088Y-0019956D02*
X0002319D01*
X0003946Y-0019990D02*
X0002270D01*
X0003824Y-0020025D02*
X0002221D01*
X0003722Y-0020059D02*
X0002172D01*
X0003626Y-0020094D02*
X0002122D01*
X0003540Y-0020129D02*
X0002073D01*
X0003459Y-0020164D02*
X0002024D01*
X0003383Y-0020198D02*
X0001982D01*
X0003315Y-0020233D02*
X0001952D01*
X0003247Y-0020268D02*
X0001922D01*
X0003185Y-0020302D02*
X0001892D01*
X0003126Y-0020337D02*
X0001862D01*
X0003067Y-0020372D02*
X0001832D01*
X0003013Y-0020407D02*
X0001802D01*
X0002962Y-0020441D02*
X0001772D01*
X0002911Y-0020476D02*
X0001742D01*
X0002862Y-0020511D02*
X0001712D01*
X0002817Y-0020545D02*
X0001682D01*
X0002773Y-0020580D02*
X0001652D01*
X0002729Y-0020615D02*
X0001622D01*
X0002687Y-0020650D02*
X0001593D01*
X0002647Y-0020684D02*
X0001563D01*
X0002608Y-0020719D02*
X0001532D01*
X0002569Y-0020754D02*
X0001502D01*
X0002532Y-0020788D02*
X0001472D01*
X0002498Y-0020823D02*
X0001443D01*
X0002463Y-0020857D02*
X0001413D01*
X0002428Y-0020892D02*
X0001390D01*
X0002395Y-0020927D02*
X0001371D01*
X0002365Y-0020962D02*
X0001352D01*
X0002334Y-0020996D02*
X0001333D01*
X0002303Y-0021031D02*
X0001314D01*
X0002273Y-0021066D02*
X0001296D01*
X0002245Y-0021100D02*
X0001277D01*
X0002218Y-0021135D02*
X0001258D01*
X0002191Y-0021170D02*
X0001239D01*
X0002164Y-0021205D02*
X0001220D01*
X0002138Y-0021239D02*
X0001202D01*
X0002114Y-0021274D02*
X0001183D01*
X0002091Y-0021309D02*
X0001164D01*
X0002067Y-0021343D02*
X0001145D01*
X0002043Y-0021378D02*
X0001126D01*
X0002020Y-0021413D02*
X0001107D01*
X0002000Y-0021447D02*
X0001089D01*
X0001979Y-0021482D02*
X0001070D01*
X0001958Y-0021517D02*
X0001051D01*
X0001938Y-0021552D02*
X0001032D01*
X0001917Y-0021586D02*
X0001013D01*
X0001899Y-0021621D02*
X0000994D01*
X0001881Y-0021656D02*
X0000976D01*
X0001864Y-0021690D02*
X0000963D01*
X0001846Y-0021725D02*
X0000952D01*
X0001828Y-0021760D02*
X0000942D01*
X0001812Y-0021794D02*
X0000931D01*
X0001797Y-0021829D02*
X0000920D01*
X0001781Y-0021864D02*
X0000910D01*
X0001766Y-0021898D02*
X0000900D01*
X0001751Y-0021933D02*
X0000889D01*
X0001736Y-0021968D02*
X0000878D01*
X0001724Y-0022002D02*
X0000868D01*
X0001711Y-0022037D02*
X0000857D01*
X0001699Y-0022072D02*
X0000847D01*
X0001686Y-0022107D02*
X0000836D01*
X0001674Y-0022141D02*
X0000826D01*
X0001662Y-0022176D02*
X0000815D01*
X0001652Y-0022211D02*
X0000805D01*
X0001642Y-0022245D02*
X0000794D01*
X0001631Y-0022280D02*
X0000783D01*
X0001621Y-0022315D02*
X0000773D01*
X0001611Y-0022350D02*
X0000763D01*
X0001602Y-0022384D02*
X0000752D01*
X0001594Y-0022419D02*
X0000741D01*
X0001587Y-0022454D02*
X0000731D01*
X0001578Y-0022488D02*
X0000720D01*
X0001570Y-0022523D02*
X0000710D01*
X0001563Y-0022557D02*
X0000699D01*
X0001556Y-0022593D02*
X0000689D01*
X0001550Y-0022627D02*
X0000687D01*
X0001544Y-0022662D02*
X0000686D01*
X0001539Y-0022696D02*
X0000684D01*
X0001533Y-0022731D02*
X0000683D01*
X0001528Y-0022766D02*
X0000681D01*
X0001523Y-0022800D02*
X0000680D01*
X0001520Y-0022835D02*
X0000678D01*
X0001517Y-0022870D02*
X0000677D01*
X0001513Y-0022905D02*
X0000676D01*
X0001510Y-0022939D02*
X0000674D01*
X0001507Y-0022974D02*
X0000672D01*
X0001504Y-0023009D02*
X0000671D01*
X0001503Y-0023043D02*
X0000670D01*
X0001502Y-0023078D02*
X0000668D01*
X0001501Y-0023113D02*
X0000667D01*
X0001500Y-0023148D02*
X0000665D01*
X0001499Y-0023182D02*
X0000664D01*
X0001498Y-0023217D02*
X0000662D01*
X0001498Y-0023252D02*
X0000661D01*
X0001500Y-0023286D02*
X0000659D01*
X0001501Y-0023321D02*
X0000658D01*
X0001502Y-0023356D02*
X0000656D01*
X0001504Y-0023390D02*
X0000655D01*
X0001505Y-0023425D02*
X0000654D01*
X0001507Y-0023460D02*
X0000652D01*
X0001511Y-0023494D02*
X0000651D01*
X0001514Y-0023529D02*
X0000649D01*
X0001517Y-0023564D02*
X0000648D01*
X0001520Y-0023598D02*
X0000656D01*
X0001524Y-0023633D02*
X0000664D01*
X0001528Y-0023668D02*
X0000671D01*
X0001533Y-0023703D02*
X0000679D01*
X0001539Y-0023737D02*
X0000687D01*
X0001545Y-0023772D02*
X0000694D01*
X0001551Y-0023807D02*
X0000702D01*
X0001556Y-0023841D02*
X0000709D01*
X0001563Y-0023876D02*
X0000717D01*
X0001570Y-0023911D02*
X0000725D01*
X0001579Y-0023945D02*
X0000732D01*
X0001587Y-0023980D02*
X0000740D01*
X0001594Y-0024015D02*
X0000748D01*
X0001603Y-0024050D02*
X0000755D01*
X0001611Y-0024084D02*
X0000763D01*
X0001622Y-0024119D02*
X0000770D01*
X0001632Y-0024154D02*
X0000778D01*
X0001643Y-0024188D02*
X0000786D01*
X0001653Y-0024223D02*
X0000793D01*
X0001664Y-0024258D02*
X0000801D01*
X0001675Y-0024293D02*
X0000809D01*
X0001688Y-0024327D02*
X0000816D01*
X0001701Y-0024362D02*
X0000824D01*
X0001713Y-0024396D02*
X0000831D01*
X0001726Y-0024431D02*
X0000839D01*
X0001739Y-0024466D02*
X0000847D01*
X0001754Y-0024500D02*
X0000854D01*
X0001769Y-0024535D02*
X0000862D01*
X0001785Y-0024570D02*
X0000877D01*
X0001800Y-0024605D02*
X0000893D01*
X0001815Y-0024639D02*
X0000910D01*
X0001831Y-0024674D02*
X0000927D01*
X0001849Y-0024709D02*
X0000943D01*
X0001867Y-0024743D02*
X0000960D01*
X0001885Y-0024778D02*
X0000977D01*
X0001903Y-0024813D02*
X0000993D01*
X0001921Y-0024848D02*
X0001010D01*
X0001942Y-0024882D02*
X0001027D01*
X0001963Y-0024917D02*
X0001043D01*
X0001983Y-0024952D02*
X0001060D01*
X0002004Y-0024986D02*
X0001077D01*
X0002025Y-0025021D02*
X0001093D01*
X0002048Y-0025056D02*
X0001110D01*
X0002072Y-0025091D02*
X0001127D01*
X0002096Y-0025125D02*
X0001143D01*
X0002120Y-0025160D02*
X0001160D01*
X0002144Y-0025194D02*
X0001177D01*
X0002170Y-0025229D02*
X0001193D01*
X0002197Y-0025264D02*
X0001210D01*
X0002224Y-0025298D02*
X0001227D01*
X0002251Y-0025333D02*
X0001243D01*
X0002278Y-0025368D02*
X0001260D01*
X0002309Y-0025403D02*
X0001277D01*
X0002340Y-0025437D02*
X0001293D01*
X0002371Y-0025472D02*
X0001310D01*
X0002402Y-0025507D02*
X0001326D01*
X0002435Y-0025541D02*
X0001343D01*
X0002469Y-0025576D02*
X0001372D01*
X0002504Y-0025611D02*
X0001405D01*
X0002538Y-0025646D02*
X0001438D01*
X0002574Y-0025680D02*
X0001471D01*
X0002614Y-0025715D02*
X0001504D01*
X0002653Y-0025750D02*
X0001537D01*
X0002693Y-0025784D02*
X0001570D01*
X0002734Y-0025819D02*
X0001603D01*
X0002779Y-0025854D02*
X0001636D01*
X0002823Y-0025888D02*
X0001669D01*
X0002867Y-0025923D02*
X0001702D01*
X0002917Y-0025958D02*
X0001735D01*
X0002968Y-0025993D02*
X0001768D01*
X0003019Y-0026027D02*
X0001800D01*
X0003072Y-0026062D02*
X0001833D01*
X0003130Y-0026096D02*
X0001867D01*
X0003188Y-0026131D02*
X0001900D01*
X0003250Y-0026166D02*
X0001933D01*
X0003317Y-0026201D02*
X0001965D01*
X0003385Y-0026235D02*
X0001998D01*
X0003459Y-0026270D02*
X0002031D01*
X0003539Y-0026305D02*
X0002065D01*
X0003622Y-0026339D02*
X0002098D01*
X0003717Y-0026374D02*
X0002130D01*
X0003816Y-0026409D02*
X0002176D01*
X0003936Y-0026443D02*
X0002227D01*
X0004072Y-0026478D02*
X0002278D01*
X0004238Y-0026513D02*
X0002330D01*
X0004496Y-0026548D02*
X0002381D01*
X0004645Y-0026582D02*
X0002432D01*
X0004645Y-0026617D02*
X0002483D01*
X0004645Y-0026652D02*
X0002534D01*
X0004645Y-0026686D02*
X0002585D01*
X0004645Y-0026721D02*
X0002636D01*
X0004645Y-0026756D02*
X0002687D01*
X0004645Y-0026791D02*
X0002739D01*
X0004645Y-0026825D02*
X0002790D01*
X0004645Y-0026860D02*
X0002841D01*
X0004645Y-0026894D02*
X0002892D01*
X0004645Y-0026929D02*
X0002952D01*
X0004645Y-0026964D02*
X0003050D01*
X0004645Y-0026998D02*
X0003149D01*
X0004645Y-0027033D02*
X0003247D01*
X0004645Y-0027068D02*
X0003346D01*
X0004645Y-0027103D02*
X0003444D01*
X0004645Y-0027137D02*
X0003542D01*
X0004645Y-0027172D02*
X0003641D01*
X0004645Y-0027207D02*
X0003739D01*
X0004645Y-0027241D02*
X0003837D01*
X0004645Y-0027276D02*
X0004051D01*
X0004645Y-0027311D02*
X0004280D01*
X0008093Y-0020678D02*
Y-0022781D01*
X0008058Y-0020644D02*
Y-0022569D01*
X0008024Y-0020611D02*
Y-0022410D01*
X0007989Y-0020578D02*
Y-0022275D01*
X0007954Y-0020544D02*
Y-0022166D01*
X0007920Y-0020511D02*
Y-0022061D01*
X0007885Y-0020477D02*
Y-0021974D01*
X0007850Y-0020444D02*
Y-0021889D01*
X0007815Y-0020410D02*
Y-0021812D01*
X0007781Y-0020377D02*
Y-0021739D01*
X0007746Y-0020343D02*
Y-0021667D01*
X0007711Y-0020310D02*
Y-0021604D01*
X0007677Y-0020277D02*
Y-0021542D01*
X0007642Y-0020243D02*
Y-0021481D01*
X0007607Y-0020210D02*
Y-0021427D01*
X0007572Y-0020176D02*
Y-0021372D01*
X0007538Y-0020143D02*
Y-0021318D01*
X0007503Y-0020109D02*
Y-0021270D01*
X0007469Y-0020076D02*
Y-0021223D01*
X0007434Y-0020043D02*
Y-0021175D01*
X0007399Y-0020009D02*
Y-0021130D01*
X0007365Y-0019978D02*
Y-0021088D01*
X0007330Y-0019955D02*
Y-0021046D01*
X0007295Y-0019931D02*
Y-0021004D01*
X0007260Y-0019908D02*
Y-0020966D01*
X0007226Y-0019885D02*
Y-0020929D01*
X0007191Y-0019861D02*
Y-0020892D01*
X0007156Y-0019838D02*
Y-0020855D01*
X0007122Y-0019815D02*
Y-0020820D01*
X0007087Y-0019791D02*
Y-0020788D01*
X0007052Y-0019768D02*
Y-0020755D01*
X0007017Y-0019744D02*
Y-0020722D01*
X0006983Y-0019721D02*
Y-0020691D01*
X0006948Y-0019698D02*
Y-0020662D01*
X0006913Y-0019674D02*
Y-0020633D01*
X0006879Y-0019651D02*
Y-0020604D01*
X0006844Y-0019628D02*
Y-0020576D01*
X0006809Y-0019604D02*
Y-0020549D01*
X0006774Y-0019581D02*
Y-0020524D01*
X0006740Y-0019557D02*
Y-0020499D01*
X0006705Y-0019534D02*
Y-0020474D01*
X0006670Y-0019511D02*
Y-0020448D01*
X0006636Y-0019487D02*
Y-0020426D01*
X0006601Y-0019474D02*
Y-0020404D01*
X0006567Y-0019463D02*
Y-0020381D01*
X0006532Y-0019450D02*
Y-0020359D01*
X0006497Y-0019438D02*
Y-0020337D01*
X0006462Y-0019426D02*
Y-0020317D01*
X0006428Y-0019414D02*
Y-0020298D01*
X0006393Y-0019402D02*
Y-0020280D01*
X0006358Y-0019390D02*
Y-0020260D01*
X0006324Y-0019378D02*
Y-0020241D01*
X0006289Y-0019366D02*
Y-0020224D01*
X0006254Y-0019354D02*
Y-0020207D01*
X0006219Y-0019341D02*
Y-0020191D01*
X0006185Y-0019330D02*
Y-0020174D01*
X0006150Y-0019317D02*
Y-0020158D01*
X0006115Y-0019305D02*
Y-0020142D01*
X0006081Y-0019293D02*
Y-0020128D01*
X0006046Y-0019281D02*
Y-0020115D01*
X0006011Y-0019269D02*
Y-0020101D01*
X0005977Y-0019257D02*
Y-0020087D01*
X0005942Y-0019244D02*
Y-0020074D01*
X0005907Y-0019233D02*
Y-0020061D01*
X0005872Y-0019220D02*
Y-0020050D01*
X0005838Y-0019208D02*
Y-0020039D01*
X0005803Y-0019196D02*
Y-0020028D01*
X0005769Y-0019184D02*
Y-0020017D01*
X0005734Y-0019175D02*
Y-0020006D01*
X0005699Y-0019172D02*
Y-0019996D01*
X0005664Y-0019169D02*
Y-0019988D01*
X0005630Y-0019165D02*
Y-0019979D01*
X0005595Y-0019162D02*
Y-0019970D01*
X0005560Y-0019159D02*
Y-0019962D01*
X0005526Y-0019156D02*
Y-0019953D01*
X0005491Y-0019153D02*
Y-0019946D01*
X0005456Y-0019150D02*
Y-0019940D01*
X0005422Y-0019146D02*
Y-0019933D01*
X0005387Y-0019143D02*
Y-0019927D01*
X0005352Y-0019140D02*
Y-0019921D01*
X0005317Y-0019137D02*
Y-0019915D01*
X0005283Y-0019133D02*
Y-0019910D01*
X0005248Y-0019130D02*
Y-0019906D01*
X0005213Y-0019127D02*
Y-0019902D01*
X0005179Y-0019124D02*
Y-0019897D01*
X0005144Y-0019120D02*
Y-0019893D01*
X0005109Y-0019117D02*
Y-0019889D01*
X0005074Y-0019114D02*
Y-0019886D01*
X0005040Y-0019111D02*
Y-0019884D01*
X0005005Y-0019108D02*
Y-0019882D01*
X0004970Y-0019105D02*
Y-0019881D01*
X0004936Y-0019101D02*
Y-0019879D01*
X0004901Y-0019098D02*
Y-0019877D01*
X0004867Y-0019095D02*
Y-0019875D01*
X0004831Y-0019092D02*
Y-0019876D01*
X0004797Y-0019089D02*
Y-0019876D01*
X0004762Y-0019085D02*
Y-0019876D01*
X0004728Y-0019082D02*
Y-0019877D01*
X0004693Y-0019086D02*
Y-0019877D01*
X0004624Y-0019096D02*
Y-0019880D01*
X0004589Y-0019102D02*
Y-0019883D01*
X0004554Y-0019107D02*
Y-0019886D01*
X0004519Y-0019112D02*
Y-0019889D01*
X0004485Y-0019117D02*
Y-0019892D01*
X0004450Y-0019122D02*
Y-0019895D01*
X0004415Y-0019127D02*
Y-0019899D01*
X0004381Y-0019132D02*
Y-0019904D01*
X0004346Y-0019137D02*
Y-0019909D01*
X0004311Y-0019143D02*
Y-0019914D01*
X0004276Y-0019148D02*
Y-0019919D01*
X0004242Y-0019153D02*
Y-0019924D01*
X0004207Y-0019157D02*
Y-0019929D01*
X0004172Y-0019163D02*
Y-0019937D01*
X0004138Y-0019168D02*
Y-0019944D01*
X0004103Y-0019173D02*
Y-0019952D01*
X0004069Y-0019178D02*
Y-0019960D01*
X0004034Y-0019183D02*
Y-0019968D01*
X0003999Y-0019188D02*
Y-0019975D01*
X0003964Y-0019193D02*
Y-0019985D01*
X0003930Y-0019198D02*
Y-0019995D01*
X0003895Y-0019204D02*
Y-0020005D01*
X0003860Y-0019209D02*
Y-0020015D01*
X0003826Y-0019214D02*
Y-0020024D01*
X0003791Y-0019223D02*
Y-0020035D01*
X0003756Y-0019236D02*
Y-0020047D01*
X0003721Y-0019250D02*
Y-0020060D01*
X0003687Y-0019263D02*
Y-0020072D01*
X0003652Y-0019276D02*
Y-0020085D01*
X0003617Y-0019289D02*
Y-0020097D01*
X0003583Y-0019302D02*
Y-0020111D01*
X0003548Y-0019315D02*
Y-0020126D01*
X0003513Y-0019328D02*
Y-0020141D01*
X0003479Y-0019342D02*
Y-0020156D01*
X0003444Y-0019355D02*
Y-0020170D01*
X0003409Y-0019368D02*
Y-0020185D01*
X0003374Y-0019381D02*
Y-0020203D01*
X0003340Y-0019394D02*
Y-0020220D01*
X0003305Y-0019407D02*
Y-0020238D01*
X0003270Y-0019421D02*
Y-0020256D01*
X0003236Y-0019434D02*
Y-0020274D01*
X0003201Y-0019447D02*
Y-0020293D01*
X0003166Y-0019460D02*
Y-0020313D01*
X0003131Y-0019474D02*
Y-0020334D01*
X0003097Y-0019487D02*
Y-0020354D01*
X0003062Y-0019500D02*
Y-0020375D01*
X0003028Y-0019513D02*
Y-0020396D01*
X0002993Y-0019526D02*
Y-0020420D01*
X0002958Y-0019539D02*
Y-0020444D01*
X0002924Y-0019553D02*
Y-0020468D01*
X0002889Y-0019566D02*
Y-0020492D01*
X0002854Y-0019579D02*
Y-0020517D01*
X0002819Y-0019603D02*
Y-0020544D01*
X0002785Y-0019628D02*
Y-0020571D01*
X0002750Y-0019652D02*
Y-0020598D01*
X0002715Y-0019677D02*
Y-0020625D01*
X0002681Y-0019701D02*
Y-0020655D01*
X0002646Y-0019726D02*
Y-0020685D01*
X0002611Y-0019750D02*
Y-0020716D01*
X0002576Y-0019774D02*
Y-0020747D01*
X0002542Y-0019799D02*
Y-0020778D01*
X0002507Y-0019823D02*
Y-0020813D01*
X0002472Y-0019848D02*
Y-0020848D01*
X0002438Y-0019872D02*
Y-0020883D01*
X0002403Y-0019896D02*
Y-0020918D01*
X0002369Y-0019921D02*
Y-0020957D01*
X0002333Y-0019946D02*
Y-0020997D01*
X0002299Y-0019970D02*
Y-0021036D01*
X0002264Y-0019994D02*
Y-0021076D01*
X0002230Y-0020019D02*
Y-0021120D01*
X0002195Y-0020043D02*
Y-0021165D01*
X0002160Y-0020068D02*
Y-0021210D01*
X0002126Y-0020092D02*
Y-0021257D01*
X0002091Y-0020117D02*
Y-0021308D01*
X0002056Y-0020141D02*
Y-0021359D01*
X0002021Y-0020165D02*
Y-0021411D01*
X0001987Y-0020193D02*
Y-0021469D01*
X0001952Y-0020233D02*
Y-0021527D01*
X0001917Y-0020273D02*
Y-0021586D01*
X0001883Y-0020313D02*
Y-0021654D01*
X0001848Y-0020354D02*
Y-0021721D01*
X0001813Y-0020394D02*
Y-0021792D01*
X0001778Y-0020434D02*
Y-0021870D01*
X0001744Y-0020474D02*
Y-0021949D01*
X0001709Y-0020514D02*
Y-0022043D01*
X0001674Y-0020554D02*
Y-0022139D01*
X0001640Y-0020594D02*
Y-0022252D01*
X0001605Y-0020635D02*
Y-0022373D01*
X0001570Y-0020675D02*
Y-0022524D01*
X0001536Y-0020715D02*
Y-0022717D01*
X0001501Y-0020756D02*
Y-0023111D01*
X0007228Y-0019886D02*
X0005082D01*
X0007280Y-0019921D02*
X0005352D01*
X0007331Y-0019956D02*
X0005535D01*
X0007380Y-0019990D02*
X0005675D01*
X0007415Y-0020025D02*
X0005794D01*
X0007452Y-0020059D02*
X0005902D01*
X0007487Y-0020094D02*
X0005994D01*
X0007524Y-0020129D02*
X0006082D01*
X0007559Y-0020164D02*
X0006162D01*
X0007595Y-0020198D02*
X0006235D01*
X0007631Y-0020233D02*
X0006308D01*
X0007667Y-0020268D02*
X0006372D01*
X0007704Y-0020302D02*
X0006435D01*
X0007739Y-0020337D02*
X0006498D01*
X0007776Y-0020372D02*
X0006552D01*
X0007811Y-0020407D02*
X0006606D01*
X0007847Y-0020441D02*
X0006660D01*
X0007883Y-0020476D02*
X0006708D01*
X0007919Y-0020511D02*
X0006756D01*
X0007956Y-0020545D02*
X0006804D01*
X0007991Y-0020580D02*
X0006849D01*
X0008028Y-0020615D02*
X0006891D01*
X0008063Y-0020650D02*
X0006933D01*
X0008100Y-0020684D02*
X0006975D01*
X0008125Y-0020719D02*
X0007014D01*
X0008146Y-0020754D02*
X0007050D01*
X0008166Y-0020788D02*
X0007087D01*
X0008187Y-0020823D02*
X0007124D01*
X0008207Y-0020857D02*
X0007159D01*
X0008227Y-0020892D02*
X0007191D01*
X0008248Y-0020927D02*
X0007224D01*
X0008268Y-0020962D02*
X0007256D01*
X0008289Y-0020996D02*
X0007289D01*
X0008309Y-0021031D02*
X0007317D01*
X0008330Y-0021066D02*
X0007346D01*
X0008350Y-0021100D02*
X0007374D01*
X0008370Y-0021135D02*
X0007403D01*
X0008391Y-0021170D02*
X0007430D01*
X0008411Y-0021205D02*
X0007455D01*
X0008432Y-0021239D02*
X0007480D01*
X0008452Y-0021274D02*
X0007506D01*
X0008472Y-0021309D02*
X0007531D01*
X0008493Y-0021343D02*
X0007554D01*
X0008513Y-0021378D02*
X0007576D01*
X0008534Y-0021413D02*
X0007598D01*
X0008554Y-0021447D02*
X0007620D01*
X0008575Y-0021482D02*
X0007643D01*
X0008595Y-0021517D02*
X0007663D01*
X0008616Y-0021552D02*
X0007682D01*
X0008636Y-0021586D02*
X0007701D01*
X0008654Y-0021621D02*
X0007720D01*
X0008664Y-0021656D02*
X0007740D01*
X0008675Y-0021690D02*
X0007757D01*
X0008686Y-0021725D02*
X0007774D01*
X0008697Y-0021760D02*
X0007791D01*
X0008707Y-0021794D02*
X0007807D01*
X0008718Y-0021829D02*
X0007824D01*
X0008729Y-0021864D02*
X0007840D01*
X0008740Y-0021898D02*
X0007854D01*
X0008751Y-0021933D02*
X0007868D01*
X0008761Y-0021968D02*
X0007882D01*
X0008772Y-0022002D02*
X0007896D01*
X0008783Y-0022037D02*
X0007910D01*
X0008794Y-0022072D02*
X0007923D01*
X0008805Y-0022107D02*
X0007935D01*
X0008815Y-0022141D02*
X0007946D01*
X0008826Y-0022176D02*
X0007957D01*
X0008837Y-0022211D02*
X0007969D01*
X0008848Y-0022245D02*
X0007980D01*
X0008859Y-0022280D02*
X0007990D01*
X0008869Y-0022315D02*
X0007999D01*
X0008880Y-0022350D02*
X0008008D01*
X0008891Y-0022384D02*
X0008017D01*
X0008902Y-0022419D02*
X0008026D01*
X0008907Y-0022454D02*
X0008035D01*
X0008909Y-0022488D02*
X0008042D01*
X0008912Y-0022523D02*
X0008049D01*
X0008914Y-0022557D02*
X0008056D01*
X0008917Y-0022593D02*
X0008063D01*
X0008919Y-0022627D02*
X0008070D01*
X-0002571Y-0024242D02*
X-0003528D01*
X-0004622D02*
X-0005576D01*
X-0000061Y-0024276D02*
X-0000978D01*
X-0002587D02*
X-0003543D01*
X-0004607D02*
X-0005560D01*
X-0000054Y-0024311D02*
X-0000972D01*
X-0002602D02*
X-0003558D01*
X-0004592D02*
X-0005544D01*
X-0000048Y-0024346D02*
X-0000965D01*
X-0002618D02*
X-0003574D01*
X-0004577D02*
X-0005529D01*
X-0000041Y-0024380D02*
X-0000959D01*
X-0002633D02*
X-0003589D01*
X-0004562D02*
X-0005513D01*
X-0000034Y-0024415D02*
X-0000952D01*
X-0002649D02*
X-0003604D01*
X-0004547D02*
X-0005498D01*
X-0000028Y-0024450D02*
X-0000945D01*
X-0002665D02*
X-0003619D01*
X-0004532D02*
X-0005483D01*
X-0000021Y-0024485D02*
X-0000939D01*
X-0002680D02*
X-0003634D01*
X-0004517D02*
X-0005467D01*
X-0000014Y-0024519D02*
X-0000932D01*
X-0002696D02*
X-0003649D01*
X-0004502D02*
X-0005452D01*
X-0000007Y-0024554D02*
X-0000926D01*
X-0002711D02*
X-0003664D01*
X-0004487D02*
X-0005436D01*
X-0000001Y-0024589D02*
X-0000919D01*
X-0002727D02*
X-0003679D01*
X-0004472D02*
X-0005420D01*
X0000005Y-0024623D02*
X-0000912D01*
X-0002743D02*
X-0003694D01*
X-0004457D02*
X-0005405D01*
X0000012Y-0024658D02*
X-0000906D01*
X-0002758D02*
X-0003709D01*
X-0004442D02*
X-0005389D01*
X0000019Y-0024693D02*
X-0000899D01*
X-0002774D02*
X-0003724D01*
X-0004427D02*
X-0005374D01*
X0000025Y-0024727D02*
X-0000893D01*
X-0002789D02*
X-0003739D01*
X-0004412D02*
X-0005358D01*
X0000032Y-0024762D02*
X-0000886D01*
X-0002805D02*
X-0003754D01*
X-0004397D02*
X-0005343D01*
X0000039Y-0024797D02*
X-0000880D01*
X-0002820D02*
X-0003769D01*
X-0004382D02*
X-0005327D01*
X0000045Y-0024831D02*
X-0000873D01*
X-0002836D02*
X-0003785D01*
X-0004367D02*
X-0005312D01*
X0000052Y-0024866D02*
X-0000866D01*
X-0002852D02*
X-0003800D01*
X-0004352D02*
X-0005296D01*
X0000059Y-0024901D02*
X-0000859D01*
X-0002867D02*
X-0003815D01*
X-0004337D02*
X-0005281D01*
X0000065Y-0024935D02*
X-0000853D01*
X-0002883D02*
X-0003830D01*
X-0004322D02*
X-0005265D01*
X0000072Y-0024970D02*
X-0000846D01*
X-0002898D02*
X-0003845D01*
X-0004307D02*
X-0005250D01*
X0000078Y-0025005D02*
X-0000840D01*
X-0002914D02*
X-0003860D01*
X-0004292D02*
X-0005234D01*
X0000085Y-0025040D02*
X-0000833D01*
X-0002930D02*
X-0003875D01*
X-0004277D02*
X-0005219D01*
X0000092Y-0025074D02*
X-0000827D01*
X-0002945D02*
X-0003890D01*
X-0004262D02*
X-0005203D01*
X0000098Y-0025109D02*
X-0000820D01*
X-0002961D02*
X-0003905D01*
X-0004247D02*
X-0005187D01*
X0000105Y-0025144D02*
X-0000813D01*
X-0002976D02*
X-0003920D01*
X-0004232D02*
X-0005172D01*
X0000112Y-0025178D02*
X-0000807D01*
X-0002992D02*
X-0003935D01*
X-0004217D02*
X-0005156D01*
X0000119Y-0025213D02*
X-0000800D01*
X-0003007D02*
X-0003950D01*
X-0004202D02*
X-0005141D01*
X0000125Y-0025248D02*
X-0000794D01*
X-0003023D02*
X-0003965D01*
X-0004187D02*
X-0005126D01*
X0000132Y-0025282D02*
X-0000787D01*
X-0003039D02*
X-0003980D01*
X-0004172D02*
X-0005110D01*
X0000139Y-0025317D02*
X-0000780D01*
X-0003054D02*
X-0003995D01*
X-0004157D02*
X-0005094D01*
X0000145Y-0025352D02*
X-0000774D01*
X-0003070D02*
X-0004011D01*
X-0004142D02*
X-0005079D01*
X0000152Y-0025387D02*
X-0000767D01*
X-0003085D02*
X-0004026D01*
X-0004127D02*
X-0005063D01*
X0000158Y-0025421D02*
X-0000761D01*
X-0003101D02*
X-0004041D01*
X-0004111D02*
X-0005048D01*
X0000165Y-0025456D02*
X-0000754D01*
X-0003117D02*
X-0004056D01*
X-0004096D02*
X-0005032D01*
X0000172Y-0025491D02*
X-0000748D01*
X-0003132D02*
X-0004071D01*
X-0004081D02*
X-0005017D01*
X0000178Y-0025525D02*
X-0000741D01*
X-0003148D02*
X-0005001D01*
X0000185Y-0025560D02*
X-0000734D01*
X-0003163D02*
X-0004986D01*
X0000192Y-0025595D02*
X-0000728D01*
X-0003179D02*
X-0004970D01*
X0000198Y-0025630D02*
X-0000721D01*
X-0003194D02*
X-0004955D01*
X0000205Y-0025664D02*
X-0000715D01*
X-0003210D02*
X-0004939D01*
X0000212Y-0025699D02*
X-0000708D01*
X-0003226D02*
X-0004924D01*
X0000219Y-0025733D02*
X-0000701D01*
X-0003241D02*
X-0004908D01*
X0000225Y-0025768D02*
X-0000695D01*
X-0003257D02*
X-0004893D01*
X0000231Y-0025803D02*
X-0000688D01*
X-0003272D02*
X-0004877D01*
X0000238Y-0025837D02*
X-0000681D01*
X-0003288D02*
X-0004861D01*
X0000245Y-0025872D02*
X-0000675D01*
X-0003304D02*
X-0004846D01*
X0000252Y-0025907D02*
X-0000668D01*
X-0003319D02*
X-0004830D01*
X0000258Y-0025942D02*
X-0000662D01*
X-0003335D02*
X-0004815D01*
X0000265Y-0025976D02*
X-0000655D01*
X-0003350D02*
X-0004800D01*
X0000272Y-0026011D02*
X-0000648D01*
X-0003366D02*
X-0004784D01*
X0000278Y-0026046D02*
X-0000642D01*
X-0003381D02*
X-0004769D01*
X0000285Y-0026080D02*
X-0000635D01*
X-0003397D02*
X-0004753D01*
X0000292Y-0026115D02*
X-0000629D01*
X-0003413D02*
X-0004737D01*
X0000298Y-0026150D02*
X-0000622D01*
X-0003428D02*
X-0004722D01*
X0000305Y-0026185D02*
X-0000615D01*
X-0003444D02*
X-0004706D01*
X0000311Y-0026219D02*
X-0000609D01*
X-0003459D02*
X-0004691D01*
X0000318Y-0026254D02*
X-0000602D01*
X-0003475D02*
X-0004675D01*
X0000325Y-0026289D02*
X-0000596D01*
X-0003491D02*
X-0004660D01*
X0000331Y-0026323D02*
X-0000589D01*
X-0003506D02*
X-0004644D01*
X0000338Y-0026358D02*
X-0000583D01*
X-0003522D02*
X-0004629D01*
X0000345Y-0026393D02*
X-0000576D01*
X-0003537D02*
X-0004613D01*
X0000352Y-0026428D02*
X-0000569D01*
X-0003553D02*
X-0004598D01*
X0000358Y-0026462D02*
X-0000563D01*
X-0003569D02*
X-0004582D01*
X0000365Y-0026497D02*
X-0000556D01*
X-0003584D02*
X-0004567D01*
X0000372Y-0026531D02*
X-0000550D01*
X-0003600D02*
X-0004551D01*
X0000378Y-0026566D02*
X-0000543D01*
X-0003615D02*
X-0004535D01*
X0000385Y-0026601D02*
X-0000536D01*
X-0003631D02*
X-0004520D01*
X0000391Y-0026635D02*
X-0000530D01*
X-0003646D02*
X-0004504D01*
X0000398Y-0026670D02*
X-0000523D01*
X-0003662D02*
X-0004489D01*
X0000405Y-0026705D02*
X-0000517D01*
X-0003678D02*
X-0004473D01*
X0000411Y-0026740D02*
X-0000510D01*
X-0003693D02*
X-0004458D01*
X0000418Y-0026774D02*
X-0000504D01*
X-0003709D02*
X-0004443D01*
X0000425Y-0026809D02*
X-0000497D01*
X-0003724D02*
X-0004427D01*
X0000431Y-0026844D02*
X-0000490D01*
X-0003740D02*
X-0004411D01*
X0000438Y-0026878D02*
X-0000483D01*
X-0003756D02*
X-0004396D01*
X0000445Y-0026913D02*
X-0000477D01*
X-0003771D02*
X-0004380D01*
X0000452Y-0026948D02*
X-0000470D01*
X-0003787D02*
X-0004365D01*
X0000458Y-0026983D02*
X-0000464D01*
X-0003802D02*
X-0004349D01*
X0000465Y-0027017D02*
X-0000457D01*
X-0003818D02*
X-0004334D01*
X0000471Y-0027052D02*
X-0000451D01*
X-0003833D02*
X-0004318D01*
X0000478Y-0027087D02*
X-0000444D01*
X-0003849D02*
X-0004303D01*
X0000485Y-0027121D02*
X-0000437D01*
X-0003865D02*
X-0004287D01*
X0000491Y-0027156D02*
X-0000431D01*
X-0003880D02*
X-0004272D01*
X0000498Y-0027191D02*
X-0000424D01*
X-0003896D02*
X-0004256D01*
X0000505Y-0027225D02*
X-0000418D01*
X-0003911D02*
X-0004241D01*
X-0004067Y-0027572D02*
X-0004085D01*
X-0007014Y-0018717D02*
X-0008654Y-0027261D01*
X-0007732D02*
X-0008654D01*
X-0006692Y-0021794D02*
X-0007732Y-0027261D01*
X-0006671Y-0021794D02*
X-0006692D01*
X-0006671D02*
X-0004076Y-0027593D01*
X-0001472Y-0021794D02*
X-0004076Y-0027593D01*
X-0001450Y-0021794D02*
X-0001472D01*
X-0001450D02*
X-0000411Y-0027261D01*
X0000512D02*
X-0000411D01*
X-0001128Y-0018717D02*
X0000512Y-0027261D01*
X-0001128Y-0018717D02*
X-0004076Y-0025503D01*
X-0007014Y-0018717D02*
X-0004076Y-0025503D01*
X0000491Y-0027152D02*
Y-0027261D01*
X0000456Y-0026971D02*
Y-0027261D01*
X0000421Y-0026791D02*
Y-0027261D01*
X0000387Y-0026610D02*
Y-0027261D01*
X0000352Y-0026429D02*
Y-0027261D01*
X0000317Y-0026248D02*
Y-0027261D01*
X0000283Y-0026067D02*
Y-0027261D01*
X0000248Y-0025887D02*
Y-0027261D01*
X0000213Y-0025706D02*
Y-0027261D01*
X0000178Y-0025525D02*
Y-0027261D01*
X0000144Y-0025344D02*
Y-0027261D01*
X0000109Y-0025164D02*
Y-0027261D01*
X0000074Y-0024983D02*
Y-0027261D01*
X0000040Y-0024802D02*
Y-0027261D01*
X0000005Y-0024621D02*
Y-0027261D01*
X-0000030Y-0024441D02*
Y-0027261D01*
X-0000064Y-0024260D02*
Y-0027261D01*
X-0000099Y-0024079D02*
Y-0027261D01*
X-0000133Y-0023898D02*
Y-0027261D01*
X-0000168Y-0023718D02*
Y-0027261D01*
X-0000203Y-0023537D02*
Y-0027261D01*
X-0000237Y-0023356D02*
Y-0027261D01*
X-0000272Y-0023176D02*
Y-0027261D01*
X-0000307Y-0022994D02*
Y-0027261D01*
X-0000342Y-0022814D02*
Y-0027261D01*
X-0000376Y-0022633D02*
Y-0027261D01*
X-0000411Y-0022452D02*
Y-0027260D01*
X-0000446Y-0022272D02*
Y-0027078D01*
X-0000480Y-0022091D02*
Y-0026895D01*
X-0000515Y-0021910D02*
Y-0026713D01*
X-0000550Y-0021730D02*
Y-0026530D01*
X-0000585Y-0021549D02*
Y-0026348D01*
X-0000619Y-0021368D02*
Y-0026165D01*
X-0000654Y-0021187D02*
Y-0025983D01*
X-0000689Y-0021006D02*
Y-0025800D01*
X-0000723Y-0020826D02*
Y-0025618D01*
X-0000758Y-0020645D02*
Y-0025435D01*
X-0000793Y-0020464D02*
Y-0025253D01*
X-0000828Y-0020283D02*
Y-0025070D01*
X-0000862Y-0020103D02*
Y-0024888D01*
X-0000897Y-0019922D02*
Y-0024706D01*
X-0000931Y-0019741D02*
Y-0024523D01*
X-0000966Y-0019560D02*
Y-0024340D01*
X-0001001Y-0019380D02*
Y-0024158D01*
X-0001035Y-0019199D02*
Y-0023975D01*
X-0001070Y-0019018D02*
Y-0023793D01*
X-0001105Y-0018837D02*
Y-0023610D01*
X-0001140Y-0018743D02*
Y-0023428D01*
X-0001174Y-0018822D02*
Y-0023245D01*
X-0001209Y-0018902D02*
Y-0023063D01*
X-0001244Y-0018982D02*
Y-0022880D01*
X-0001278Y-0019062D02*
Y-0022698D01*
X-0001313Y-0019142D02*
Y-0022515D01*
X-0001348Y-0019222D02*
Y-0022333D01*
X-0001383Y-0019302D02*
Y-0022150D01*
X-0001417Y-0019382D02*
Y-0021968D01*
X-0001452Y-0019461D02*
Y-0021794D01*
X-0001487Y-0019541D02*
Y-0021826D01*
X-0001521Y-0019621D02*
Y-0021904D01*
X-0001556Y-0019701D02*
Y-0021981D01*
X-0001591Y-0019781D02*
Y-0022058D01*
X-0001625Y-0019861D02*
Y-0022135D01*
X-0001660Y-0019941D02*
Y-0022213D01*
X-0001695Y-0020020D02*
Y-0022290D01*
X-0001730Y-0020100D02*
Y-0022367D01*
X-0001764Y-0020180D02*
Y-0022444D01*
X-0001799Y-0020260D02*
Y-0022522D01*
X-0001833Y-0020340D02*
Y-0022599D01*
X-0001868Y-0020420D02*
Y-0022676D01*
X-0001903Y-0020500D02*
Y-0022753D01*
X-0001938Y-0020580D02*
Y-0022831D01*
X-0001972Y-0020659D02*
Y-0022908D01*
X-0002007Y-0020739D02*
Y-0022985D01*
X-0002042Y-0020819D02*
Y-0023062D01*
X-0002076Y-0020899D02*
Y-0023140D01*
X-0002111Y-0020979D02*
Y-0023217D01*
X-0002146Y-0021059D02*
Y-0023294D01*
X-0002180Y-0021139D02*
Y-0023371D01*
X-0002215Y-0021219D02*
Y-0023448D01*
X-0002250Y-0021298D02*
Y-0023526D01*
X-0002285Y-0021378D02*
Y-0023603D01*
X-0002319Y-0021458D02*
Y-0023680D01*
X-0002354Y-0021538D02*
Y-0023757D01*
X-0002389Y-0021618D02*
Y-0023835D01*
X-0002423Y-0021698D02*
Y-0023912D01*
X-0002458Y-0021778D02*
Y-0023989D01*
X-0002493Y-0021858D02*
Y-0024067D01*
X-0002528Y-0021937D02*
Y-0024144D01*
X-0002562Y-0022017D02*
Y-0024221D01*
X-0002597Y-0022097D02*
Y-0024298D01*
X-0002631Y-0022177D02*
Y-0024376D01*
X-0002666Y-0022257D02*
Y-0024453D01*
X-0002701Y-0022337D02*
Y-0024530D01*
X-0002735Y-0022417D02*
Y-0024607D01*
X-0002770Y-0022496D02*
Y-0024685D01*
X-0002805Y-0022576D02*
Y-0024762D01*
X-0002840Y-0022656D02*
Y-0024839D01*
X-0002874Y-0022736D02*
Y-0024917D01*
X-0002909Y-0022816D02*
Y-0024994D01*
X-0002944Y-0022896D02*
Y-0025071D01*
X-0002978Y-0022976D02*
Y-0025148D01*
X-0003013Y-0023056D02*
Y-0025226D01*
X-0003048Y-0023135D02*
Y-0025303D01*
X-0003083Y-0023215D02*
Y-0025380D01*
X-0003117Y-0023295D02*
Y-0025457D01*
X-0003152Y-0023375D02*
Y-0025535D01*
X-0003187Y-0023455D02*
Y-0025612D01*
X-0003221Y-0023535D02*
Y-0025689D01*
X-0003256Y-0023615D02*
Y-0025767D01*
X-0003291Y-0023695D02*
Y-0025844D01*
X-0003326Y-0023774D02*
Y-0025921D01*
X-0003360Y-0023854D02*
Y-0025998D01*
X-0003395Y-0023934D02*
Y-0026075D01*
X-0003430Y-0024014D02*
Y-0026153D01*
X-0003464Y-0024094D02*
Y-0026230D01*
X-0003499Y-0024174D02*
Y-0026307D01*
X-0003533Y-0024254D02*
Y-0026384D01*
X-0003568Y-0024334D02*
Y-0026462D01*
X-0003603Y-0024413D02*
Y-0026539D01*
X-0003638Y-0024493D02*
Y-0026616D01*
X-0003672Y-0024573D02*
Y-0026693D01*
X-0003707Y-0024653D02*
Y-0026771D01*
X-0003742Y-0024733D02*
Y-0026848D01*
X-0003776Y-0024813D02*
Y-0026925D01*
X-0003811Y-0024893D02*
Y-0027002D01*
X-0003846Y-0024972D02*
Y-0027080D01*
X-0003881Y-0025052D02*
Y-0027157D01*
X-0003915Y-0025132D02*
Y-0027234D01*
X-0003950Y-0025212D02*
Y-0027311D01*
X-0003985Y-0025292D02*
Y-0027389D01*
X-0004019Y-0025372D02*
Y-0027466D01*
X-0004054Y-0025452D02*
Y-0027543D01*
X-0004089Y-0025474D02*
Y-0027565D01*
X-0004123Y-0025394D02*
Y-0027487D01*
X-0004158Y-0025314D02*
Y-0027410D01*
X-0004193Y-0025233D02*
Y-0027332D01*
X-0004228Y-0025154D02*
Y-0027255D01*
X-0004262Y-0025073D02*
Y-0027177D01*
X-0004297Y-0024993D02*
Y-0027100D01*
X-0004331Y-0024913D02*
Y-0027022D01*
X-0004366Y-0024833D02*
Y-0026944D01*
X-0004401Y-0024753D02*
Y-0026867D01*
X-0004436Y-0024672D02*
Y-0026789D01*
X-0004470Y-0024593D02*
Y-0026712D01*
X-0004505Y-0024512D02*
Y-0026634D01*
X-0004540Y-0024432D02*
Y-0026557D01*
X-0004574Y-0024352D02*
Y-0026479D01*
X-0004609Y-0024272D02*
Y-0026402D01*
X-0004644Y-0024192D02*
Y-0026324D01*
X-0004678Y-0024111D02*
Y-0026246D01*
X-0004713Y-0024031D02*
Y-0026169D01*
X-0004748Y-0023951D02*
Y-0026091D01*
X-0004783Y-0023871D02*
Y-0026014D01*
X-0004817Y-0023791D02*
Y-0025937D01*
X-0004852Y-0023711D02*
Y-0025859D01*
X-0004887Y-0023631D02*
Y-0025781D01*
X-0004921Y-0023550D02*
Y-0025704D01*
X-0004956Y-0023470D02*
Y-0025626D01*
X-0004991Y-0023390D02*
Y-0025549D01*
X-0005026Y-0023310D02*
Y-0025471D01*
X-0005060Y-0023230D02*
Y-0025394D01*
X-0005095Y-0023150D02*
Y-0025316D01*
X-0005130Y-0023070D02*
Y-0025239D01*
X-0005164Y-0022989D02*
Y-0025161D01*
X-0005199Y-0022909D02*
Y-0025083D01*
X-0005233Y-0022829D02*
Y-0025006D01*
X-0005269Y-0022749D02*
Y-0024928D01*
X-0005303Y-0022669D02*
Y-0024851D01*
X-0005338Y-0022589D02*
Y-0024773D01*
X-0005372Y-0022509D02*
Y-0024696D01*
X-0005407Y-0022428D02*
Y-0024618D01*
X-0005442Y-0022348D02*
Y-0024541D01*
X-0005476Y-0022268D02*
Y-0024463D01*
X-0005511Y-0022188D02*
Y-0024386D01*
X-0005546Y-0022108D02*
Y-0024308D01*
X-0005581Y-0022028D02*
Y-0024231D01*
X-0005615Y-0021948D02*
Y-0024153D01*
X-0005650Y-0021867D02*
Y-0024076D01*
X-0005685Y-0021787D02*
Y-0023998D01*
X-0005719Y-0021707D02*
Y-0023920D01*
X-0005754Y-0021627D02*
Y-0023843D01*
X-0005789Y-0021547D02*
Y-0023765D01*
X-0005824Y-0021467D02*
Y-0023688D01*
X-0005858Y-0021387D02*
Y-0023610D01*
X-0005893Y-0021306D02*
Y-0023533D01*
X-0005928Y-0021226D02*
Y-0023455D01*
X-0005962Y-0021146D02*
Y-0023378D01*
X-0005997Y-0021066D02*
Y-0023300D01*
X-0006031Y-0020986D02*
Y-0023222D01*
X-0006066Y-0020906D02*
Y-0023145D01*
X-0006101Y-0020826D02*
Y-0023067D01*
X-0006136Y-0020745D02*
Y-0022990D01*
X-0006170Y-0020665D02*
Y-0022913D01*
X-0006205Y-0020585D02*
Y-0022835D01*
X-0006240Y-0020505D02*
Y-0022757D01*
X-0006274Y-0020425D02*
Y-0022680D01*
X-0006309Y-0020344D02*
Y-0022602D01*
X-0006344Y-0020265D02*
Y-0022525D01*
X-0006379Y-0020184D02*
Y-0022447D01*
X-0006413Y-0020104D02*
Y-0022370D01*
X-0006448Y-0020024D02*
Y-0022292D01*
X-0006483Y-0019944D02*
Y-0022215D01*
X-0006517Y-0019864D02*
Y-0022137D01*
X-0006552Y-0019783D02*
Y-0022059D01*
X-0006587Y-0019704D02*
Y-0021982D01*
X-0006621Y-0019623D02*
Y-0021904D01*
X-0006656Y-0019543D02*
Y-0021827D01*
X-0006691Y-0019463D02*
Y-0021794D01*
X-0006726Y-0019383D02*
Y-0021971D01*
X-0006760Y-0019303D02*
Y-0022153D01*
X-0006795Y-0019222D02*
Y-0022335D01*
X-0006830Y-0019142D02*
Y-0022518D01*
X-0006864Y-0019062D02*
Y-0022700D01*
X-0006899Y-0018982D02*
Y-0022882D01*
X-0006934Y-0018902D02*
Y-0023065D01*
X-0006969Y-0018822D02*
Y-0023247D01*
X-0007003Y-0018742D02*
Y-0023430D01*
X-0007038Y-0018840D02*
Y-0023612D01*
X-0007072Y-0019021D02*
Y-0023794D01*
X-0007107Y-0019202D02*
Y-0023976D01*
X-0007142Y-0019382D02*
Y-0024159D01*
X-0007176Y-0019563D02*
Y-0024341D01*
X-0007211Y-0019744D02*
Y-0024524D01*
X-0007246Y-0019925D02*
Y-0024706D01*
X-0007281Y-0020106D02*
Y-0024888D01*
X-0007315Y-0020286D02*
Y-0025071D01*
X-0007350Y-0020467D02*
Y-0025253D01*
X-0007385Y-0020648D02*
Y-0025435D01*
X-0007419Y-0020828D02*
Y-0025618D01*
X-0007454Y-0021009D02*
Y-0025800D01*
X-0007489Y-0021190D02*
Y-0025982D01*
X-0007524Y-0021371D02*
Y-0026165D01*
X-0007558Y-0021552D02*
Y-0026347D01*
X-0007593Y-0021732D02*
Y-0026530D01*
X-0007628Y-0021913D02*
Y-0026712D01*
X-0007662Y-0022094D02*
Y-0026894D01*
X-0007697Y-0022274D02*
Y-0027076D01*
X-0007731Y-0022455D02*
Y-0027259D01*
X-0007767Y-0022636D02*
Y-0027261D01*
X-0007801Y-0022817D02*
Y-0027261D01*
X-0007836Y-0022998D02*
Y-0027261D01*
X-0007870Y-0023178D02*
Y-0027261D01*
X-0007905Y-0023359D02*
Y-0027261D01*
X-0007940Y-0023540D02*
Y-0027261D01*
X-0007974Y-0023720D02*
Y-0027261D01*
X-0008009Y-0023901D02*
Y-0027261D01*
X-0008044Y-0024082D02*
Y-0027261D01*
X-0008079Y-0024263D02*
Y-0027261D01*
X-0008113Y-0024444D02*
Y-0027261D01*
X-0008148Y-0024624D02*
Y-0027261D01*
X-0008183Y-0024805D02*
Y-0027261D01*
X-0008217Y-0024986D02*
Y-0027261D01*
X-0008252Y-0025167D02*
Y-0027261D01*
X-0008287Y-0025347D02*
Y-0027261D01*
X-0008322Y-0025528D02*
Y-0027261D01*
X-0008356Y-0025709D02*
Y-0027261D01*
X-0008391Y-0025889D02*
Y-0027261D01*
X-0008426Y-0026070D02*
Y-0027261D01*
X-0008460Y-0026251D02*
Y-0027261D01*
X-0008495Y-0026432D02*
Y-0027261D01*
X-0008530Y-0026613D02*
Y-0027261D01*
X-0008564Y-0026793D02*
Y-0027261D01*
X-0008599Y-0026974D02*
Y-0027261D01*
X-0008634Y-0027155D02*
Y-0027261D01*
X-0006995Y-0018760D02*
X-0007022D01*
X-0006980Y-0018794D02*
X-0007029D01*
X-0006965Y-0018829D02*
X-0007036D01*
X-0006950Y-0018864D02*
X-0007042D01*
X-0006935Y-0018898D02*
X-0007049D01*
X-0006920Y-0018933D02*
X-0007056D01*
X-0006905Y-0018968D02*
X-0007062D01*
X-0006890Y-0019003D02*
X-0007069D01*
X-0006875Y-0019037D02*
X-0007076D01*
X-0006860Y-0019072D02*
X-0007082D01*
X-0006845Y-0019107D02*
X-0007089D01*
X-0006830Y-0019141D02*
X-0007096D01*
X-0006815Y-0019176D02*
X-0007102D01*
X-0006800Y-0019211D02*
X-0007109D01*
X-0006785Y-0019246D02*
X-0007115D01*
X-0006770Y-0019280D02*
X-0007122D01*
X-0006755Y-0019315D02*
X-0007129D01*
X-0006740Y-0019350D02*
X-0007135D01*
X-0006725Y-0019384D02*
X-0007142D01*
X-0006710Y-0019419D02*
X-0007149D01*
X-0006695Y-0019454D02*
X-0007156D01*
X-0006680Y-0019489D02*
X-0007162D01*
X-0006665Y-0019523D02*
X-0007169D01*
X-0006650Y-0019558D02*
X-0007176D01*
X-0006635Y-0019593D02*
X-0007182D01*
X-0006620Y-0019627D02*
X-0007189D01*
X-0006605Y-0019662D02*
X-0007195D01*
X-0006590Y-0019696D02*
X-0007202D01*
X-0006575Y-0019731D02*
X-0007209D01*
X-0006559Y-0019766D02*
X-0007215D01*
X-0006544Y-0019801D02*
X-0007222D01*
X-0006530Y-0019835D02*
X-0007229D01*
X-0006515Y-0019870D02*
X-0007235D01*
X-0006500Y-0019905D02*
X-0007242D01*
X-0006485Y-0019939D02*
X-0007249D01*
X-0006470Y-0019974D02*
X-0007256D01*
X-0006454Y-0020009D02*
X-0007262D01*
X-0006439Y-0020044D02*
X-0007269D01*
X-0006424Y-0020078D02*
X-0007275D01*
X-0006409Y-0020113D02*
X-0007282D01*
X-0006394Y-0020148D02*
X-0007289D01*
X-0006380Y-0020182D02*
X-0007295D01*
X-0006365Y-0020217D02*
X-0007302D01*
X-0006349Y-0020252D02*
X-0007309D01*
X-0006334Y-0020286D02*
X-0007315D01*
X-0006319Y-0020321D02*
X-0007322D01*
X-0006304Y-0020356D02*
X-0007329D01*
X-0006289Y-0020391D02*
X-0007335D01*
X-0006274Y-0020425D02*
X-0007342D01*
X-0006259Y-0020460D02*
X-0007349D01*
X-0006244Y-0020494D02*
X-0007355D01*
X-0006229Y-0020529D02*
X-0007362D01*
X-0006214Y-0020564D02*
X-0007369D01*
X-0006199Y-0020599D02*
X-0007375D01*
X-0006184Y-0020633D02*
X-0007382D01*
X-0006169Y-0020668D02*
X-0007389D01*
X-0006154Y-0020703D02*
X-0007395D01*
X-0006139Y-0020737D02*
X-0007402D01*
X-0006124Y-0020772D02*
X-0007409D01*
X-0006109Y-0020807D02*
X-0007415D01*
X-0006094Y-0020841D02*
X-0007422D01*
X-0006079Y-0020876D02*
X-0007429D01*
X-0006064Y-0020911D02*
X-0007435D01*
X-0006049Y-0020946D02*
X-0007442D01*
X-0006034Y-0020980D02*
X-0007448D01*
X-0006019Y-0021015D02*
X-0007455D01*
X-0006004Y-0021050D02*
X-0007462D01*
X-0005989Y-0021084D02*
X-0007469D01*
X-0005974Y-0021119D02*
X-0007475D01*
X-0005959Y-0021154D02*
X-0007482D01*
X-0005944Y-0021189D02*
X-0007489D01*
X-0005929Y-0021223D02*
X-0007495D01*
X-0005914Y-0021258D02*
X-0007502D01*
X-0005899Y-0021293D02*
X-0007508D01*
X-0005884Y-0021327D02*
X-0007515D01*
X-0005869Y-0021362D02*
X-0007522D01*
X-0005854Y-0021396D02*
X-0007528D01*
X-0005839Y-0021431D02*
X-0007535D01*
X-0005824Y-0021466D02*
X-0007542D01*
X-0005809Y-0021501D02*
X-0007548D01*
X-0005794Y-0021535D02*
X-0007555D01*
X-0005779Y-0021570D02*
X-0007562D01*
X-0005764Y-0021605D02*
X-0007569D01*
X-0005748Y-0021639D02*
X-0007575D01*
X-0005733Y-0021674D02*
X-0007582D01*
X-0005719Y-0021709D02*
X-0007588D01*
X-0005704Y-0021744D02*
X-0007595D01*
X-0005689Y-0021778D02*
X-0007602D01*
X-0006696Y-0021813D02*
X-0007608D01*
X-0006702Y-0021848D02*
X-0007615D01*
X-0006709Y-0021882D02*
X-0007622D01*
X-0006715Y-0021917D02*
X-0007628D01*
X-0006722Y-0021952D02*
X-0007635D01*
X-0006728Y-0021987D02*
X-0007642D01*
X-0006735Y-0022021D02*
X-0007648D01*
X-0006742Y-0022056D02*
X-0007655D01*
X-0006748Y-0022091D02*
X-0007662D01*
X-0006755Y-0022125D02*
X-0007668D01*
X-0006761Y-0022160D02*
X-0007675D01*
X-0006768Y-0022194D02*
X-0007681D01*
X-0006775Y-0022229D02*
X-0007688D01*
X-0006781Y-0022264D02*
X-0007695D01*
X-0006788Y-0022299D02*
X-0007702D01*
X-0006794Y-0022333D02*
X-0007708D01*
X-0006801Y-0022368D02*
X-0007715D01*
X-0006808Y-0022403D02*
X-0007722D01*
X-0006814Y-0022437D02*
X-0007728D01*
X-0006821Y-0022472D02*
X-0007735D01*
X-0006828Y-0022507D02*
X-0007742D01*
X-0006834Y-0022542D02*
X-0007748D01*
X-0006841Y-0022576D02*
X-0007755D01*
X-0006847Y-0022611D02*
X-0007761D01*
X-0006854Y-0022646D02*
X-0007768D01*
X-0006861Y-0022680D02*
X-0007775D01*
X-0006867Y-0022715D02*
X-0007781D01*
X-0006874Y-0022750D02*
X-0007788D01*
X-0006880Y-0022784D02*
X-0007795D01*
X-0006887Y-0022819D02*
X-0007802D01*
X-0006894Y-0022854D02*
X-0007808D01*
X-0006900Y-0022889D02*
X-0007815D01*
X-0006907Y-0022923D02*
X-0007822D01*
X-0006913Y-0022958D02*
X-0007828D01*
X-0006920Y-0022993D02*
X-0007835D01*
X-0006926Y-0023027D02*
X-0007841D01*
X-0006933Y-0023062D02*
X-0007848D01*
X-0006940Y-0023097D02*
X-0007855D01*
X-0006946Y-0023131D02*
X-0007861D01*
X-0006953Y-0023166D02*
X-0007868D01*
X-0006959Y-0023201D02*
X-0007875D01*
X-0006966Y-0023235D02*
X-0007881D01*
X-0006973Y-0023270D02*
X-0007888D01*
X-0006979Y-0023305D02*
X-0007895D01*
X-0006986Y-0023339D02*
X-0007902D01*
X-0006993Y-0023374D02*
X-0007908D01*
X-0006999Y-0023409D02*
X-0007915D01*
X-0007006Y-0023444D02*
X-0007921D01*
X-0007012Y-0023478D02*
X-0007928D01*
X-0007019Y-0023513D02*
X-0007935D01*
X-0007026Y-0023548D02*
X-0007941D01*
X-0007032Y-0023582D02*
X-0007948D01*
X-0007039Y-0023617D02*
X-0007955D01*
X-0007045Y-0023652D02*
X-0007961D01*
X-0007052Y-0023687D02*
X-0007968D01*
X-0007059Y-0023721D02*
X-0007975D01*
X-0007065Y-0023756D02*
X-0007981D01*
X-0007072Y-0023791D02*
X-0007988D01*
X-0007078Y-0023825D02*
X-0007994D01*
X-0007085Y-0023860D02*
X-0008001D01*
X-0007092Y-0023894D02*
X-0008008D01*
X-0007098Y-0023930D02*
X-0008015D01*
X-0007105Y-0023964D02*
X-0008021D01*
X-0007111Y-0023999D02*
X-0008028D01*
X-0007118Y-0024033D02*
X-0008035D01*
X-0007124Y-0024068D02*
X-0008041D01*
X-0007131Y-0024103D02*
X-0008048D01*
X-0007138Y-0024137D02*
X-0008055D01*
X-0007144Y-0024172D02*
X-0008061D01*
X-0007151Y-0024207D02*
X-0008068D01*
X-0007157Y-0024242D02*
X-0008074D01*
X-0007164Y-0024276D02*
X-0008081D01*
X-0007171Y-0024311D02*
X-0008088D01*
X-0007178Y-0024346D02*
X-0008094D01*
X-0007184Y-0024380D02*
X-0008101D01*
X-0007191Y-0024415D02*
X-0008108D01*
X-0007197Y-0024450D02*
X-0008115D01*
X-0007204Y-0024485D02*
X-0008121D01*
X-0007210Y-0024519D02*
X-0008128D01*
X-0007217Y-0024554D02*
X-0008135D01*
X-0007224Y-0024589D02*
X-0008141D01*
X-0007230Y-0024623D02*
X-0008148D01*
X-0007237Y-0024658D02*
X-0008154D01*
X-0007243Y-0024693D02*
X-0008161D01*
X-0007250Y-0024727D02*
X-0008168D01*
X-0007257Y-0024762D02*
X-0008174D01*
X-0007263Y-0024797D02*
X-0008181D01*
X-0007270Y-0024831D02*
X-0008188D01*
X-0007276Y-0024866D02*
X-0008194D01*
X-0007283Y-0024901D02*
X-0008201D01*
X-0007290Y-0024935D02*
X-0008208D01*
X-0007296Y-0024970D02*
X-0008215D01*
X-0007303Y-0025005D02*
X-0008221D01*
X-0007309Y-0025040D02*
X-0008228D01*
X-0007316Y-0025074D02*
X-0008234D01*
X-0007322Y-0025109D02*
X-0008241D01*
X-0007329Y-0025144D02*
X-0008248D01*
X-0007336Y-0025178D02*
X-0008254D01*
X-0007343Y-0025213D02*
X-0008261D01*
X-0007349Y-0025248D02*
X-0008268D01*
X-0007356Y-0025282D02*
X-0008274D01*
X-0007362Y-0025317D02*
X-0008281D01*
X-0007369Y-0025352D02*
X-0008288D01*
X-0007376Y-0025387D02*
X-0008294D01*
X-0007382Y-0025421D02*
X-0008301D01*
X-0007389Y-0025456D02*
X-0008307D01*
X-0007395Y-0025491D02*
X-0008314D01*
X-0007402Y-0025525D02*
X-0008321D01*
X-0007408Y-0025560D02*
X-0008328D01*
X-0007415Y-0025595D02*
X-0008334D01*
X-0007422Y-0025630D02*
X-0008341D01*
X-0007428Y-0025664D02*
X-0008348D01*
X-0007435Y-0025699D02*
X-0008354D01*
X-0007441Y-0025733D02*
X-0008361D01*
X-0007448Y-0025768D02*
X-0008368D01*
X-0007455Y-0025803D02*
X-0008374D01*
X-0007461Y-0025837D02*
X-0008381D01*
X-0007468Y-0025872D02*
X-0008387D01*
X-0007474Y-0025907D02*
X-0008394D01*
X-0007481Y-0025942D02*
X-0008401D01*
X-0007488Y-0025976D02*
X-0008407D01*
X-0007494Y-0026011D02*
X-0008414D01*
X-0007501Y-0026046D02*
X-0008421D01*
X-0007507Y-0026080D02*
X-0008428D01*
X-0007514Y-0026115D02*
X-0008434D01*
X-0007520Y-0026150D02*
X-0008441D01*
X-0007527Y-0026185D02*
X-0008448D01*
X-0007534Y-0026219D02*
X-0008454D01*
X-0007541Y-0026254D02*
X-0008461D01*
X-0007547Y-0026289D02*
X-0008467D01*
X-0007554Y-0026323D02*
X-0008474D01*
X-0007560Y-0026358D02*
X-0008481D01*
X-0007567Y-0026393D02*
X-0008487D01*
X-0007574Y-0026428D02*
X-0008494D01*
X-0007580Y-0026462D02*
X-0008501D01*
X-0007587Y-0026497D02*
X-0008507D01*
X-0007593Y-0026531D02*
X-0008514D01*
X-0007600Y-0026566D02*
X-0008521D01*
X-0007606Y-0026601D02*
X-0008528D01*
X-0007613Y-0026635D02*
X-0008534D01*
X-0007620Y-0026670D02*
X-0008541D01*
X-0007626Y-0026705D02*
X-0008547D01*
X-0007633Y-0026740D02*
X-0008554D01*
X-0007639Y-0026774D02*
X-0008561D01*
X-0007646Y-0026809D02*
X-0008567D01*
X-0007653Y-0026844D02*
X-0008574D01*
X-0007659Y-0026878D02*
X-0008581D01*
X-0007666Y-0026913D02*
X-0008587D01*
X-0007672Y-0026948D02*
X-0008594D01*
X-0007679Y-0026983D02*
X-0008601D01*
X-0007686Y-0027017D02*
X-0008607D01*
X-0007692Y-0027052D02*
X-0008614D01*
X-0007699Y-0027087D02*
X-0008620D01*
X-0007706Y-0027121D02*
X-0008627D01*
X-0007712Y-0027156D02*
X-0008634D01*
X-0007719Y-0027191D02*
X-0008641D01*
X-0007725Y-0027225D02*
X-0008647D01*
X-0003927Y-0027260D02*
X-0004225D01*
X-0003943Y-0027295D02*
X-0004209D01*
X-0003958Y-0027330D02*
X-0004194D01*
X-0003974Y-0027364D02*
X-0004178D01*
X-0003989Y-0027399D02*
X-0004163D01*
X-0004005Y-0027433D02*
X-0004147D01*
X-0004020Y-0027468D02*
X-0004132D01*
X-0004036Y-0027503D02*
X-0004117D01*
X-0004052Y-0027538D02*
X-0004101D01*
X-0001120Y-0018760D02*
X-0001147D01*
X-0001113Y-0018794D02*
X-0001162D01*
X-0001106Y-0018829D02*
X-0001177D01*
X-0001100Y-0018864D02*
X-0001192D01*
X-0001093Y-0018898D02*
X-0001207D01*
X-0001087Y-0018933D02*
X-0001222D01*
X-0001080Y-0018968D02*
X-0001237D01*
X-0001073Y-0019003D02*
X-0001252D01*
X-0001067Y-0019037D02*
X-0001268D01*
X-0001060Y-0019072D02*
X-0001283D01*
X-0001053Y-0019107D02*
X-0001298D01*
X-0001046Y-0019141D02*
X-0001313D01*
X-0001040Y-0019176D02*
X-0001328D01*
X-0001033Y-0019211D02*
X-0001343D01*
X-0001027Y-0019246D02*
X-0001358D01*
X-0001020Y-0019280D02*
X-0001373D01*
X-0001013Y-0019315D02*
X-0001388D01*
X-0001007Y-0019350D02*
X-0001403D01*
X-0001000Y-0019384D02*
X-0001418D01*
X-0000993Y-0019419D02*
X-0001433D01*
X-0000987Y-0019454D02*
X-0001448D01*
X-0000980Y-0019489D02*
X-0001463D01*
X-0000973Y-0019523D02*
X-0001479D01*
X-0000967Y-0019558D02*
X-0001494D01*
X-0000960Y-0019593D02*
X-0001509D01*
X-0000953Y-0019627D02*
X-0001524D01*
X-0000947Y-0019662D02*
X-0001539D01*
X-0000940Y-0019696D02*
X-0001554D01*
X-0000933Y-0019731D02*
X-0001569D01*
X-0000927Y-0019766D02*
X-0001584D01*
X-0000920Y-0019801D02*
X-0001599D01*
X-0000913Y-0019835D02*
X-0001614D01*
X-0000907Y-0019870D02*
X-0001629D01*
X-0000900Y-0019905D02*
X-0001644D01*
X-0000893Y-0019939D02*
X-0001659D01*
X-0000887Y-0019974D02*
X-0001674D01*
X-0000880Y-0020009D02*
X-0001690D01*
X-0000873Y-0020044D02*
X-0001705D01*
X-0000867Y-0020078D02*
X-0001720D01*
X-0000860Y-0020113D02*
X-0001735D01*
X-0000854Y-0020148D02*
X-0001750D01*
X-0000847Y-0020182D02*
X-0001765D01*
X-0000840Y-0020217D02*
X-0001780D01*
X-0000833Y-0020252D02*
X-0001795D01*
X-0000827Y-0020286D02*
X-0001810D01*
X-0000820Y-0020321D02*
X-0001825D01*
X-0000813Y-0020356D02*
X-0001840D01*
X-0000807Y-0020391D02*
X-0001856D01*
X-0000800Y-0020425D02*
X-0001870D01*
X-0000793Y-0020460D02*
X-0001885D01*
X-0000787Y-0020494D02*
X-0001900D01*
X-0000780Y-0020529D02*
X-0001916D01*
X-0000774Y-0020564D02*
X-0001931D01*
X-0000767Y-0020599D02*
X-0001946D01*
X-0000760Y-0020633D02*
X-0001961D01*
X-0000754Y-0020668D02*
X-0001976D01*
X-0000747Y-0020703D02*
X-0001991D01*
X-0000740Y-0020737D02*
X-0002006D01*
X-0000733Y-0020772D02*
X-0002021D01*
X-0000727Y-0020807D02*
X-0002036D01*
X-0000720Y-0020841D02*
X-0002051D01*
X-0000713Y-0020876D02*
X-0002067D01*
X-0000707Y-0020911D02*
X-0002081D01*
X-0000700Y-0020946D02*
X-0002096D01*
X-0000694Y-0020980D02*
X-0002111D01*
X-0000687Y-0021015D02*
X-0002127D01*
X-0000680Y-0021050D02*
X-0002142D01*
X-0000674Y-0021084D02*
X-0002157D01*
X-0000667Y-0021119D02*
X-0002172D01*
X-0000660Y-0021154D02*
X-0002187D01*
X-0000654Y-0021189D02*
X-0002202D01*
X-0000647Y-0021223D02*
X-0002217D01*
X-0000640Y-0021258D02*
X-0002232D01*
X-0000634Y-0021293D02*
X-0002247D01*
X-0000627Y-0021327D02*
X-0002262D01*
X-0000620Y-0021362D02*
X-0002277D01*
X-0000614Y-0021396D02*
X-0002293D01*
X-0000607Y-0021431D02*
X-0002307D01*
X-0000600Y-0021466D02*
X-0002322D01*
X-0000594Y-0021501D02*
X-0002338D01*
X-0000587Y-0021535D02*
X-0002353D01*
X-0000580Y-0021570D02*
X-0002368D01*
X-0000574Y-0021605D02*
X-0002383D01*
X-0000567Y-0021639D02*
X-0002398D01*
X-0000560Y-0021674D02*
X-0002413D01*
X-0000554Y-0021709D02*
X-0002428D01*
X-0000547Y-0021744D02*
X-0002443D01*
X-0000541Y-0021778D02*
X-0002458D01*
X-0000534Y-0021813D02*
X-0001446D01*
X-0001481D02*
X-0002473D01*
X-0005674D02*
X-0006662D01*
X-0000527Y-0021848D02*
X-0001440D01*
X-0001496D02*
X-0002488D01*
X-0005659D02*
X-0006647D01*
X-0000520Y-0021882D02*
X-0001433D01*
X-0001512D02*
X-0002504D01*
X-0005643D02*
X-0006631D01*
X-0000514Y-0021917D02*
X-0001427D01*
X-0001527D02*
X-0002519D01*
X-0005628D02*
X-0006616D01*
X-0000507Y-0021952D02*
X-0001420D01*
X-0001543D02*
X-0002533D01*
X-0005613D02*
X-0006600D01*
X-0000500Y-0021987D02*
X-0001414D01*
X-0001559D02*
X-0002549D01*
X-0005598D02*
X-0006585D01*
X-0000494Y-0022021D02*
X-0001407D01*
X-0001574D02*
X-0002564D01*
X-0005583D02*
X-0006569D01*
X-0000487Y-0022056D02*
X-0001400D01*
X-0001590D02*
X-0002579D01*
X-0005569D02*
X-0006554D01*
X-0000480Y-0022091D02*
X-0001394D01*
X-0001605D02*
X-0002594D01*
X-0005554D02*
X-0006538D01*
X-0000474Y-0022125D02*
X-0001387D01*
X-0001621D02*
X-0002609D01*
X-0005538D02*
X-0006522D01*
X-0000467Y-0022160D02*
X-0001381D01*
X-0001637D02*
X-0002624D01*
X-0005523D02*
X-0006507D01*
X-0000461Y-0022194D02*
X-0001374D01*
X-0001652D02*
X-0002639D01*
X-0005508D02*
X-0006492D01*
X-0000454Y-0022229D02*
X-0001367D01*
X-0001668D02*
X-0002654D01*
X-0005493D02*
X-0006476D01*
X-0000447Y-0022264D02*
X-0001361D01*
X-0001683D02*
X-0002669D01*
X-0005478D02*
X-0006461D01*
X-0000441Y-0022299D02*
X-0001354D01*
X-0001699D02*
X-0002684D01*
X-0005463D02*
X-0006445D01*
X-0000434Y-0022333D02*
X-0001348D01*
X-0001714D02*
X-0002699D01*
X-0005448D02*
X-0006430D01*
X-0000427Y-0022368D02*
X-0001341D01*
X-0001730D02*
X-0002715D01*
X-0005433D02*
X-0006414D01*
X-0000420Y-0022403D02*
X-0001335D01*
X-0001746D02*
X-0002730D01*
X-0005418D02*
X-0006398D01*
X-0000414Y-0022437D02*
X-0001328D01*
X-0001761D02*
X-0002744D01*
X-0005403D02*
X-0006383D01*
X-0000407Y-0022472D02*
X-0001321D01*
X-0001777D02*
X-0002759D01*
X-0005388D02*
X-0006367D01*
X-0000400Y-0022507D02*
X-0001315D01*
X-0001792D02*
X-0002775D01*
X-0005373D02*
X-0006352D01*
X-0000394Y-0022542D02*
X-0001308D01*
X-0001808D02*
X-0002790D01*
X-0005358D02*
X-0006336D01*
X-0000387Y-0022576D02*
X-0001302D01*
X-0001823D02*
X-0002805D01*
X-0005343D02*
X-0006321D01*
X-0000381Y-0022611D02*
X-0001295D01*
X-0001839D02*
X-0002820D01*
X-0005328D02*
X-0006305D01*
X-0000374Y-0022646D02*
X-0001288D01*
X-0001855D02*
X-0002835D01*
X-0005313D02*
X-0006290D01*
X-0000367Y-0022680D02*
X-0001282D01*
X-0001870D02*
X-0002850D01*
X-0005298D02*
X-0006274D01*
X-0000361Y-0022715D02*
X-0001275D01*
X-0001886D02*
X-0002865D01*
X-0005283D02*
X-0006259D01*
X-0000354Y-0022750D02*
X-0001269D01*
X-0001901D02*
X-0002880D01*
X-0005268D02*
X-0006243D01*
X-0000347Y-0022784D02*
X-0001262D01*
X-0001917D02*
X-0002895D01*
X-0005253D02*
X-0006228D01*
X-0000341Y-0022819D02*
X-0001256D01*
X-0001932D02*
X-0002910D01*
X-0005238D02*
X-0006212D01*
X-0000334Y-0022854D02*
X-0001249D01*
X-0001948D02*
X-0002926D01*
X-0005223D02*
X-0006196D01*
X-0000327Y-0022889D02*
X-0001242D01*
X-0001964D02*
X-0002941D01*
X-0005208D02*
X-0006181D01*
X-0000320Y-0022923D02*
X-0001235D01*
X-0001979D02*
X-0002956D01*
X-0005193D02*
X-0006166D01*
X-0000314Y-0022958D02*
X-0001229D01*
X-0001995D02*
X-0002970D01*
X-0005178D02*
X-0006150D01*
X-0000307Y-0022993D02*
X-0001222D01*
X-0002010D02*
X-0002986D01*
X-0005163D02*
X-0006135D01*
X-0000301Y-0023027D02*
X-0001216D01*
X-0002026D02*
X-0003001D01*
X-0005148D02*
X-0006119D01*
X-0000294Y-0023062D02*
X-0001209D01*
X-0002041D02*
X-0003016D01*
X-0005133D02*
X-0006104D01*
X-0000287Y-0023097D02*
X-0001203D01*
X-0002057D02*
X-0003031D01*
X-0005118D02*
X-0006088D01*
X-0000281Y-0023131D02*
X-0001196D01*
X-0002073D02*
X-0003046D01*
X-0005103D02*
X-0006072D01*
X-0000274Y-0023166D02*
X-0001189D01*
X-0002088D02*
X-0003061D01*
X-0005088D02*
X-0006057D01*
X-0000267Y-0023201D02*
X-0001183D01*
X-0002104D02*
X-0003076D01*
X-0005073D02*
X-0006041D01*
X-0000261Y-0023235D02*
X-0001176D01*
X-0002119D02*
X-0003091D01*
X-0005058D02*
X-0006026D01*
X-0000254Y-0023270D02*
X-0001170D01*
X-0002135D02*
X-0003106D01*
X-0005043D02*
X-0006010D01*
X-0000247Y-0023305D02*
X-0001163D01*
X-0002150D02*
X-0003121D01*
X-0005028D02*
X-0005995D01*
X-0000241Y-0023339D02*
X-0001156D01*
X-0002166D02*
X-0003136D01*
X-0005013D02*
X-0005979D01*
X-0000234Y-0023374D02*
X-0001150D01*
X-0002182D02*
X-0003152D01*
X-0004998D02*
X-0005964D01*
X-0000228Y-0023409D02*
X-0001143D01*
X-0002197D02*
X-0003167D01*
X-0004983D02*
X-0005948D01*
X-0000221Y-0023444D02*
X-0001137D01*
X-0002213D02*
X-0003181D01*
X-0004968D02*
X-0005933D01*
X-0000214Y-0023478D02*
X-0001130D01*
X-0002228D02*
X-0003197D01*
X-0004953D02*
X-0005917D01*
X-0000207Y-0023513D02*
X-0001124D01*
X-0002244D02*
X-0003212D01*
X-0004937D02*
X-0005902D01*
X-0000201Y-0023548D02*
X-0001117D01*
X-0002260D02*
X-0003227D01*
X-0004922D02*
X-0005886D01*
X-0000194Y-0023582D02*
X-0001110D01*
X-0002275D02*
X-0003242D01*
X-0004907D02*
X-0005870D01*
X-0000187Y-0023617D02*
X-0001104D01*
X-0002291D02*
X-0003257D01*
X-0004893D02*
X-0005855D01*
X-0000181Y-0023652D02*
X-0001097D01*
X-0002306D02*
X-0003272D01*
X-0004878D02*
X-0005839D01*
X-0000174Y-0023687D02*
X-0001091D01*
X-0002322D02*
X-0003287D01*
X-0004863D02*
X-0005824D01*
X-0000167Y-0023721D02*
X-0001084D01*
X-0002337D02*
X-0003302D01*
X-0004848D02*
X-0005809D01*
X-0000161Y-0023756D02*
X-0001077D01*
X-0002353D02*
X-0003317D01*
X-0004832D02*
X-0005793D01*
X-0000154Y-0023791D02*
X-0001070D01*
X-0002369D02*
X-0003332D01*
X-0004817D02*
X-0005778D01*
X-0000148Y-0023825D02*
X-0001064D01*
X-0002384D02*
X-0003347D01*
X-0004802D02*
X-0005762D01*
X-0000141Y-0023860D02*
X-0001057D01*
X-0002400D02*
X-0003363D01*
X-0004787D02*
X-0005746D01*
X-0000134Y-0023894D02*
X-0001051D01*
X-0002415D02*
X-0003378D01*
X-0004772D02*
X-0005731D01*
X-0000128Y-0023930D02*
X-0001044D01*
X-0002431D02*
X-0003393D01*
X-0004757D02*
X-0005715D01*
X-0000121Y-0023964D02*
X-0001038D01*
X-0002446D02*
X-0003408D01*
X-0004743D02*
X-0005700D01*
X-0000114Y-0023999D02*
X-0001031D01*
X-0002462D02*
X-0003423D01*
X-0004727D02*
X-0005684D01*
X-0000107Y-0024033D02*
X-0001024D01*
X-0002478D02*
X-0003438D01*
X-0004712D02*
X-0005669D01*
X-0000101Y-0024068D02*
X-0001018D01*
X-0002493D02*
X-0003453D01*
X-0004697D02*
X-0005653D01*
X-0000094Y-0024103D02*
X-0001011D01*
X-0002509D02*
X-0003468D01*
X-0004682D02*
X-0005638D01*
X-0000087Y-0024137D02*
X-0001005D01*
X-0002524D02*
X-0003483D01*
X-0004667D02*
X-0005622D01*
X-0000081Y-0024172D02*
X-0000998D01*
X-0002540D02*
X-0003498D01*
X-0004652D02*
X-0005607D01*
X-0000074Y-0024207D02*
X-0000991D01*
X-0002556D02*
X-0003513D01*
X-0004637D02*
X-0005591D01*
X-0000068Y-0024242D02*
X-0000985D01*
X-0010463Y-0019178D02*
Y-0021002D01*
X-0010498Y-0019178D02*
Y-0021052D01*
X-0010533Y-0019178D02*
Y-0021102D01*
X-0010567Y-0019178D02*
Y-0021153D01*
X-0010602Y-0019178D02*
Y-0021204D01*
X-0010637Y-0019178D02*
Y-0021254D01*
X-0010671Y-0019178D02*
Y-0021305D01*
X-0010706Y-0019178D02*
Y-0021355D01*
X-0010741Y-0019178D02*
Y-0021406D01*
X-0010776Y-0019178D02*
Y-0021456D01*
X-0010810Y-0019178D02*
Y-0021507D01*
X-0010845Y-0019178D02*
Y-0021557D01*
X-0010880Y-0019178D02*
Y-0021607D01*
X-0010914Y-0019178D02*
Y-0021658D01*
X-0010949Y-0019178D02*
Y-0021709D01*
X-0010984Y-0019178D02*
Y-0021759D01*
X-0011019Y-0019178D02*
Y-0021810D01*
X-0011053Y-0019178D02*
Y-0021860D01*
X-0011088Y-0019178D02*
Y-0021911D01*
X-0011122Y-0019178D02*
Y-0021961D01*
X-0011157Y-0019178D02*
Y-0022012D01*
X-0011192Y-0019178D02*
Y-0022062D01*
X-0011226Y-0019178D02*
Y-0022113D01*
X-0011261Y-0019178D02*
Y-0022163D01*
X-0011296Y-0019178D02*
Y-0022214D01*
X-0011331Y-0019178D02*
Y-0022265D01*
X-0011365Y-0019178D02*
Y-0022315D01*
X-0011400Y-0019178D02*
Y-0022365D01*
X-0011435Y-0019178D02*
Y-0022416D01*
X-0011469Y-0019178D02*
Y-0022467D01*
X-0011504Y-0019178D02*
Y-0022517D01*
X-0011539Y-0019178D02*
Y-0022568D01*
X-0011574Y-0019178D02*
Y-0022618D01*
X-0011608Y-0019178D02*
Y-0022669D01*
X-0011643Y-0019178D02*
Y-0022719D01*
X-0011678Y-0019178D02*
Y-0022770D01*
X-0011712Y-0019178D02*
Y-0022820D01*
X-0011747Y-0019178D02*
Y-0022870D01*
X-0011781Y-0019178D02*
Y-0022921D01*
X-0014280Y-0019178D02*
Y-0022913D01*
X-0014315Y-0019178D02*
Y-0022862D01*
X-0014349Y-0019178D02*
Y-0022812D01*
X-0014384Y-0019178D02*
Y-0022761D01*
X-0014419Y-0019178D02*
Y-0022711D01*
X-0014453Y-0019178D02*
Y-0022660D01*
X-0014488Y-0019178D02*
Y-0022609D01*
X-0014522Y-0019178D02*
Y-0022559D01*
X-0014557Y-0019178D02*
Y-0022508D01*
X-0014592Y-0019178D02*
Y-0022458D01*
X-0014627Y-0019178D02*
Y-0022407D01*
X-0014661Y-0019178D02*
Y-0022357D01*
X-0014696Y-0019178D02*
Y-0022306D01*
X-0014731Y-0019178D02*
Y-0022256D01*
X-0014765Y-0019178D02*
Y-0022205D01*
X-0014800Y-0019178D02*
Y-0022155D01*
X-0014835Y-0019178D02*
Y-0022104D01*
X-0014870Y-0019178D02*
Y-0022054D01*
X-0014904Y-0019178D02*
Y-0022003D01*
X-0014939Y-0019178D02*
Y-0021952D01*
X-0014974Y-0019178D02*
Y-0021902D01*
X-0015008Y-0019178D02*
Y-0021852D01*
X-0015043Y-0019178D02*
Y-0021801D01*
X-0015078Y-0019178D02*
Y-0021750D01*
X-0015112Y-0019178D02*
Y-0021700D01*
X-0015147Y-0019178D02*
Y-0021649D01*
X-0015182Y-0019178D02*
Y-0021599D01*
X-0015217Y-0019178D02*
Y-0021548D01*
X-0015251Y-0019178D02*
Y-0021498D01*
X-0015286Y-0019178D02*
Y-0021447D01*
X-0015320Y-0019178D02*
Y-0021397D01*
X-0015355Y-0019178D02*
Y-0021346D01*
X-0015390Y-0019178D02*
Y-0021296D01*
X-0015425Y-0019178D02*
Y-0021245D01*
X-0015459Y-0019178D02*
Y-0021194D01*
X-0015494Y-0019178D02*
Y-0021144D01*
X-0015529Y-0019178D02*
Y-0021093D01*
X-0015563Y-0019178D02*
Y-0021043D01*
X-0015598Y-0019178D02*
Y-0020993D01*
X-0015633Y-0019178D02*
Y-0020942D01*
X-0015667Y-0019178D02*
Y-0020891D01*
X-0015702Y-0019178D02*
Y-0020841D01*
X-0015737Y-0019178D02*
Y-0020790D01*
X-0015772Y-0019178D02*
Y-0020740D01*
X-0015806Y-0019178D02*
Y-0020689D01*
X-0015841Y-0019178D02*
Y-0020639D01*
X-0015876Y-0019178D02*
Y-0020588D01*
X-0015910Y-0019178D02*
Y-0020537D01*
X-0015945Y-0019178D02*
Y-0020487D01*
X-0015980Y-0019178D02*
Y-0020437D01*
X-0016015Y-0019178D02*
Y-0020386D01*
X-0016049Y-0019178D02*
Y-0020335D01*
X-0016084Y-0019178D02*
Y-0020285D01*
X-0016119Y-0019178D02*
Y-0020234D01*
X-0016153Y-0019178D02*
Y-0020184D01*
X-0016188Y-0019178D02*
Y-0020133D01*
X-0016222Y-0019178D02*
Y-0020083D01*
X-0016257Y-0019178D02*
Y-0020032D01*
X-0016292Y-0019178D02*
Y-0019981D01*
X-0016327Y-0019178D02*
Y-0019931D01*
X-0016361Y-0019178D02*
Y-0019881D01*
X-0016396Y-0019178D02*
Y-0019830D01*
X-0016431Y-0019178D02*
Y-0019780D01*
X-0016465Y-0019178D02*
Y-0019729D01*
X-0016500Y-0019178D02*
Y-0019678D01*
X-0016535Y-0019178D02*
Y-0019628D01*
X-0016570Y-0019178D02*
Y-0019578D01*
X-0016604Y-0019178D02*
Y-0019527D01*
X-0016639Y-0019178D02*
Y-0019476D01*
X-0016674Y-0019178D02*
Y-0019426D01*
X-0016708Y-0019178D02*
Y-0019375D01*
X-0016743Y-0019178D02*
Y-0019325D01*
X-0016778Y-0019178D02*
Y-0019274D01*
X-0016813Y-0019178D02*
Y-0019224D01*
X-0009220Y-0019192D02*
X-0011803D01*
X-0009244Y-0019226D02*
X-0011824D01*
X-0009268Y-0019261D02*
X-0011844D01*
X-0009292Y-0019296D02*
X-0011865D01*
X-0009316Y-0019330D02*
X-0011885D01*
X-0009339Y-0019365D02*
X-0011906D01*
X-0009363Y-0019400D02*
X-0011926D01*
X-0009387Y-0019435D02*
X-0011946D01*
X-0009411Y-0019469D02*
X-0011967D01*
X-0009435Y-0019504D02*
X-0011987D01*
X-0009459Y-0019539D02*
X-0012007D01*
X-0009482Y-0019573D02*
X-0012028D01*
X-0009506Y-0019608D02*
X-0012048D01*
X-0009530Y-0019643D02*
X-0012069D01*
X-0009554Y-0019677D02*
X-0012089D01*
X-0009578Y-0019712D02*
X-0012110D01*
X-0009602Y-0019747D02*
X-0012130D01*
X-0009625Y-0019781D02*
X-0012151D01*
X-0009649Y-0019816D02*
X-0012171D01*
X-0009673Y-0019851D02*
X-0012192D01*
X-0009697Y-0019885D02*
X-0012212D01*
X-0009721Y-0019920D02*
X-0012233D01*
X-0009744Y-0019955D02*
X-0012253D01*
X-0009769Y-0019990D02*
X-0012273D01*
X-0009792Y-0020024D02*
X-0012294D01*
X-0009816Y-0020059D02*
X-0012314D01*
X-0009840Y-0020094D02*
X-0012335D01*
X-0009864Y-0020128D02*
X-0012355D01*
X-0009887Y-0020163D02*
X-0012376D01*
X-0009911Y-0020198D02*
X-0012396D01*
X-0009935Y-0020232D02*
X-0012417D01*
X-0009959Y-0020267D02*
X-0012437D01*
X-0009983Y-0020302D02*
X-0012457D01*
X-0010007Y-0020337D02*
X-0012478D01*
X-0010030Y-0020371D02*
X-0012498D01*
X-0010054Y-0020406D02*
X-0012519D01*
X-0010078Y-0020441D02*
X-0012539D01*
X-0010102Y-0020475D02*
X-0012559D01*
X-0010126Y-0020510D02*
X-0012580D01*
X-0010150Y-0020545D02*
X-0012600D01*
X-0010173Y-0020580D02*
X-0012621D01*
X-0010197Y-0020614D02*
X-0012641D01*
X-0010221Y-0020649D02*
X-0012662D01*
X-0010245Y-0020683D02*
X-0012682D01*
X-0010269Y-0020718D02*
X-0012703D01*
X-0010293Y-0020753D02*
X-0012723D01*
X-0010317Y-0020787D02*
X-0012744D01*
X-0010340Y-0020822D02*
X-0012764D01*
X-0010364Y-0020857D02*
X-0012785D01*
X-0010388Y-0020892D02*
X-0012805D01*
X-0010412Y-0020926D02*
X-0012825D01*
X-0010435Y-0020961D02*
X-0012846D01*
X-0010459Y-0020996D02*
X-0012866D01*
X-0010483Y-0021030D02*
X-0012887D01*
X-0010507Y-0021065D02*
X-0012907D01*
X-0010531Y-0021100D02*
X-0012928D01*
X-0010555Y-0021135D02*
X-0012948D01*
X-0010578Y-0021169D02*
X-0012969D01*
X-0010602Y-0021204D02*
X-0012989D01*
X-0010626Y-0021239D02*
X-0013009D01*
X-0010620Y-0024639D02*
X-0013018D01*
X-0010595Y-0024673D02*
X-0012996D01*
X-0010571Y-0024708D02*
X-0012974D01*
X-0010547Y-0024743D02*
X-0012951D01*
X-0010523Y-0024778D02*
X-0012929D01*
X-0010499Y-0024812D02*
X-0012907D01*
X-0010475Y-0024847D02*
X-0012884D01*
X-0010451Y-0024881D02*
X-0012862D01*
X-0010427Y-0024916D02*
X-0012840D01*
X-0010403Y-0024951D02*
X-0012817D01*
X-0010379Y-0024986D02*
X-0012795D01*
X-0010355Y-0025020D02*
X-0012773D01*
X-0010331Y-0025055D02*
X-0012751D01*
X-0010307Y-0025090D02*
X-0012728D01*
X-0010283Y-0025124D02*
X-0012706D01*
X-0010259Y-0025159D02*
X-0012684D01*
X-0010235Y-0025194D02*
X-0012661D01*
X-0010211Y-0025228D02*
X-0012639D01*
X-0010187Y-0025263D02*
X-0012617D01*
X-0010163Y-0025298D02*
X-0012594D01*
X-0010139Y-0025333D02*
X-0012572D01*
X-0010115Y-0025367D02*
X-0012550D01*
X-0010091Y-0025402D02*
X-0012528D01*
X-0010067Y-0025437D02*
X-0012506D01*
X-0010043Y-0025471D02*
X-0012483D01*
X-0010019Y-0025506D02*
X-0012461D01*
X-0009995Y-0025541D02*
X-0012439D01*
X-0009971Y-0025576D02*
X-0012417D01*
X-0009947Y-0025610D02*
X-0012394D01*
X-0009923Y-0025645D02*
X-0012372D01*
X-0009899Y-0025680D02*
X-0012350D01*
X-0009875Y-0025714D02*
X-0012327D01*
X-0009851Y-0025749D02*
X-0012305D01*
X-0009827Y-0025783D02*
X-0012283D01*
X-0009803Y-0025819D02*
X-0012260D01*
X-0009779Y-0025853D02*
X-0012238D01*
X-0009755Y-0025888D02*
X-0012216D01*
X-0009731Y-0025922D02*
X-0012194D01*
X-0009707Y-0025957D02*
X-0012171D01*
X-0009683Y-0025992D02*
X-0012149D01*
X-0009659Y-0026026D02*
X-0012127D01*
X-0009635Y-0026061D02*
X-0012104D01*
X-0009611Y-0026096D02*
X-0012082D01*
X-0009587Y-0026131D02*
X-0012060D01*
X-0009563Y-0026165D02*
X-0012037D01*
X-0009539Y-0026200D02*
X-0012015D01*
X-0009515Y-0026235D02*
X-0011993D01*
X-0009491Y-0026269D02*
X-0011971D01*
X-0009467Y-0026304D02*
X-0011948D01*
X-0009443Y-0026339D02*
X-0011926D01*
X-0009419Y-0026374D02*
X-0011904D01*
X-0009394Y-0026408D02*
X-0011881D01*
X-0009370Y-0026443D02*
X-0011859D01*
X-0009346Y-0026478D02*
X-0011837D01*
X-0009322Y-0026512D02*
X-0011815D01*
X-0009298Y-0026547D02*
X-0011793D01*
X-0009274Y-0026581D02*
X-0011770D01*
X-0009250Y-0026616D02*
X-0011748D01*
X-0009226Y-0026651D02*
X-0011726D01*
X-0009202Y-0026686D02*
X-0011703D01*
X-0009178Y-0026720D02*
X-0011681D01*
X-0009154Y-0026755D02*
X-0011659D01*
X-0009130Y-0026790D02*
X-0011637D01*
X-0009106Y-0026824D02*
X-0011614D01*
X-0009082Y-0026859D02*
X-0011592D01*
X-0009058Y-0026894D02*
X-0011570D01*
X-0009034Y-0026929D02*
X-0011547D01*
X-0009010Y-0026963D02*
X-0011525D01*
X-0008986Y-0026998D02*
X-0011503D01*
X-0008962Y-0027033D02*
X-0011480D01*
X-0008938Y-0027067D02*
X-0011458D01*
X-0008914Y-0027102D02*
X-0011436D01*
X-0008890Y-0027137D02*
X-0011414D01*
X-0008866Y-0027171D02*
X-0011391D01*
X-0008842Y-0027206D02*
X-0011369D01*
X-0008818Y-0027241D02*
X-0011347D01*
X-0014868D02*
X-0017408D01*
X-0014261Y-0019178D02*
X-0016844D01*
X-0014261D02*
X-0013028Y-0021269D01*
X-0011795Y-0019178D02*
X-0013028Y-0021269D01*
X-0009211Y-0019178D02*
X-0011795D01*
X-0009211D02*
X-0011795Y-0022941D01*
X-0008804Y-0027261D01*
X-0011334D01*
X-0013028Y-0024624D02*
X-0011334Y-0027261D01*
X-0013028Y-0024624D02*
X-0014883Y-0027261D01*
X-0017423D01*
X-0014261Y-0022941D02*
X-0017423Y-0027261D01*
X-0016844Y-0019178D02*
X-0014261Y-0022941D01*
X-0008833Y-0027220D02*
Y-0027261D01*
X-0008867Y-0027169D02*
Y-0027261D01*
X-0008902Y-0027119D02*
Y-0027261D01*
X-0008937Y-0027069D02*
Y-0027261D01*
X-0008971Y-0027019D02*
Y-0027261D01*
X-0009006Y-0026969D02*
Y-0027261D01*
X-0009041Y-0026919D02*
Y-0027261D01*
X-0009076Y-0026869D02*
Y-0027261D01*
X-0009110Y-0026819D02*
Y-0027261D01*
X-0009145Y-0026769D02*
Y-0027261D01*
X-0009180Y-0026719D02*
Y-0027261D01*
X-0009214Y-0026669D02*
Y-0027261D01*
X-0009249Y-0026618D02*
Y-0027261D01*
X-0009283Y-0026568D02*
Y-0027261D01*
X-0009319Y-0026518D02*
Y-0027261D01*
X-0009353Y-0026468D02*
Y-0027261D01*
X-0009388Y-0026418D02*
Y-0027261D01*
X-0009422Y-0026368D02*
Y-0027261D01*
X-0009457Y-0026318D02*
Y-0027261D01*
X-0009492Y-0026267D02*
Y-0027261D01*
X-0009526Y-0026217D02*
Y-0027261D01*
X-0009561Y-0026167D02*
Y-0027261D01*
X-0009596Y-0026117D02*
Y-0027261D01*
X-0009631Y-0026067D02*
Y-0027261D01*
X-0009665Y-0026017D02*
Y-0027261D01*
X-0009700Y-0025967D02*
Y-0027261D01*
X-0009735Y-0025917D02*
Y-0027261D01*
X-0009769Y-0025867D02*
Y-0027261D01*
X-0009804Y-0025817D02*
Y-0027261D01*
X-0009839Y-0025767D02*
Y-0027261D01*
X-0009874Y-0025716D02*
Y-0027261D01*
X-0009908Y-0025666D02*
Y-0027261D01*
X-0009943Y-0025616D02*
Y-0027261D01*
X-0009978Y-0025566D02*
Y-0027261D01*
X-0010012Y-0025516D02*
Y-0027261D01*
X-0010047Y-0025466D02*
Y-0027261D01*
X-0010081Y-0025416D02*
Y-0027261D01*
X-0010116Y-0025365D02*
Y-0027261D01*
X-0010151Y-0025315D02*
Y-0027261D01*
X-0010186Y-0025265D02*
Y-0027261D01*
X-0010220Y-0025215D02*
Y-0027261D01*
X-0010255Y-0025165D02*
Y-0027261D01*
X-0010290Y-0025115D02*
Y-0027261D01*
X-0010324Y-0025065D02*
Y-0027261D01*
X-0010359Y-0025015D02*
Y-0027261D01*
X-0010394Y-0024965D02*
Y-0027261D01*
X-0010429Y-0024915D02*
Y-0027261D01*
X-0010463Y-0024864D02*
Y-0027261D01*
X-0010498Y-0024814D02*
Y-0027261D01*
X-0010533Y-0024764D02*
Y-0027261D01*
X-0010567Y-0024714D02*
Y-0027261D01*
X-0010602Y-0024664D02*
Y-0027261D01*
X-0010637Y-0024614D02*
Y-0027261D01*
X-0010671Y-0024564D02*
Y-0027261D01*
X-0010706Y-0024514D02*
Y-0027261D01*
X-0010741Y-0024463D02*
Y-0027261D01*
X-0010776Y-0024413D02*
Y-0027261D01*
X-0010810Y-0024363D02*
Y-0027261D01*
X-0010845Y-0024313D02*
Y-0027261D01*
X-0010880Y-0024263D02*
Y-0027261D01*
X-0010914Y-0024213D02*
Y-0027261D01*
X-0010949Y-0024163D02*
Y-0027261D01*
X-0010984Y-0024113D02*
Y-0027261D01*
X-0011019Y-0024063D02*
Y-0027261D01*
X-0011053Y-0024013D02*
Y-0027261D01*
X-0011088Y-0023962D02*
Y-0027261D01*
X-0011122Y-0023912D02*
Y-0027261D01*
X-0011157Y-0023862D02*
Y-0027261D01*
X-0011192Y-0023812D02*
Y-0027261D01*
X-0011226Y-0023762D02*
Y-0027261D01*
X-0011261Y-0023712D02*
Y-0027261D01*
X-0011296Y-0023662D02*
Y-0027261D01*
X-0011331Y-0023611D02*
Y-0027261D01*
X-0011365Y-0023561D02*
Y-0027212D01*
X-0011400Y-0023511D02*
Y-0027158D01*
X-0011435Y-0023461D02*
Y-0027104D01*
X-0011469Y-0023411D02*
Y-0027050D01*
X-0011504Y-0023361D02*
Y-0026996D01*
X-0011539Y-0023311D02*
Y-0026942D01*
X-0011574Y-0023261D02*
Y-0026888D01*
X-0011608Y-0023211D02*
Y-0026834D01*
X-0011643Y-0023161D02*
Y-0026780D01*
X-0011678Y-0023111D02*
Y-0026726D01*
X-0011712Y-0023060D02*
Y-0026672D01*
X-0011747Y-0023010D02*
Y-0026618D01*
X-0011781Y-0022960D02*
Y-0026564D01*
X-0011817Y-0019214D02*
Y-0026510D01*
X-0011851Y-0019273D02*
Y-0026456D01*
X-0011886Y-0019331D02*
Y-0026402D01*
X-0011920Y-0019391D02*
Y-0026348D01*
X-0011955Y-0019449D02*
Y-0026294D01*
X-0011990Y-0019508D02*
Y-0026240D01*
X-0012024Y-0019567D02*
Y-0026185D01*
X-0012059Y-0019626D02*
Y-0026131D01*
X-0012094Y-0019685D02*
Y-0026078D01*
X-0012129Y-0019744D02*
Y-0026024D01*
X-0012163Y-0019803D02*
Y-0025970D01*
X-0012198Y-0019861D02*
Y-0025915D01*
X-0012233Y-0019920D02*
Y-0025861D01*
X-0012267Y-0019979D02*
Y-0025807D01*
X-0012302Y-0020038D02*
Y-0025754D01*
X-0012337Y-0020097D02*
Y-0025700D01*
X-0012372Y-0020156D02*
Y-0025645D01*
X-0012406Y-0020215D02*
Y-0025591D01*
X-0012441Y-0020274D02*
Y-0025537D01*
X-0012476Y-0020333D02*
Y-0025483D01*
X-0012510Y-0020391D02*
Y-0025430D01*
X-0012545Y-0020450D02*
Y-0025375D01*
X-0012580Y-0020509D02*
Y-0025321D01*
X-0012614Y-0020568D02*
Y-0025267D01*
X-0012649Y-0020627D02*
Y-0025213D01*
X-0012684Y-0020686D02*
Y-0025159D01*
X-0012719Y-0020745D02*
Y-0025105D01*
X-0012753Y-0020804D02*
Y-0025051D01*
X-0012788Y-0020863D02*
Y-0024997D01*
X-0012822Y-0020921D02*
Y-0024943D01*
X-0012857Y-0020980D02*
Y-0024889D01*
X-0012892Y-0021039D02*
Y-0024835D01*
X-0012927Y-0021098D02*
Y-0024781D01*
X-0012961Y-0021157D02*
Y-0024727D01*
X-0012996Y-0021216D02*
Y-0024673D01*
X-0013031Y-0021263D02*
Y-0024629D01*
X-0013065Y-0021205D02*
Y-0024678D01*
X-0013100Y-0021146D02*
Y-0024728D01*
X-0013135Y-0021087D02*
Y-0024777D01*
X-0013169Y-0021028D02*
Y-0024826D01*
X-0013204Y-0020969D02*
Y-0024876D01*
X-0013239Y-0020911D02*
Y-0024925D01*
X-0013274Y-0020852D02*
Y-0024974D01*
X-0013308Y-0020793D02*
Y-0025024D01*
X-0013343Y-0020734D02*
Y-0025073D01*
X-0013378Y-0020675D02*
Y-0025122D01*
X-0013412Y-0020616D02*
Y-0025171D01*
X-0013447Y-0020557D02*
Y-0025221D01*
X-0013482Y-0020498D02*
Y-0025270D01*
X-0013517Y-0020440D02*
Y-0025319D01*
X-0013551Y-0020381D02*
Y-0025369D01*
X-0013586Y-0020322D02*
Y-0025418D01*
X-0013620Y-0020263D02*
Y-0025467D01*
X-0013655Y-0020204D02*
Y-0025517D01*
X-0013690Y-0020145D02*
Y-0025566D01*
X-0013724Y-0020087D02*
Y-0025615D01*
X-0013759Y-0020028D02*
Y-0025665D01*
X-0013794Y-0019969D02*
Y-0025714D01*
X-0013829Y-0019910D02*
Y-0025763D01*
X-0013863Y-0019851D02*
Y-0025813D01*
X-0013898Y-0019793D02*
Y-0025862D01*
X-0013933Y-0019733D02*
Y-0025911D01*
X-0013967Y-0019675D02*
Y-0025961D01*
X-0014002Y-0019616D02*
Y-0026010D01*
X-0014037Y-0019557D02*
Y-0026059D01*
X-0014072Y-0019498D02*
Y-0026108D01*
X-0014106Y-0019439D02*
Y-0026158D01*
X-0014141Y-0019380D02*
Y-0026207D01*
X-0014176Y-0019322D02*
Y-0026256D01*
X-0014210Y-0019263D02*
Y-0026306D01*
X-0014245Y-0019204D02*
Y-0026355D01*
X-0014280Y-0022967D02*
Y-0026404D01*
X-0014315Y-0023015D02*
Y-0026454D01*
X-0014349Y-0023062D02*
Y-0026503D01*
X-0014384Y-0023109D02*
Y-0026552D01*
X-0014419Y-0023157D02*
Y-0026602D01*
X-0014453Y-0023204D02*
Y-0026651D01*
X-0014488Y-0023252D02*
Y-0026700D01*
X-0014522Y-0023299D02*
Y-0026750D01*
X-0014557Y-0023346D02*
Y-0026799D01*
X-0014592Y-0023394D02*
Y-0026848D01*
X-0014627Y-0023441D02*
Y-0026898D01*
X-0014661Y-0023489D02*
Y-0026947D01*
X-0014696Y-0023536D02*
Y-0026996D01*
X-0014731Y-0023583D02*
Y-0027046D01*
X-0014765Y-0023631D02*
Y-0027095D01*
X-0014800Y-0023678D02*
Y-0027144D01*
X-0014835Y-0023726D02*
Y-0027193D01*
X-0014870Y-0023773D02*
Y-0027243D01*
X-0014904Y-0023820D02*
Y-0027261D01*
X-0014939Y-0023868D02*
Y-0027261D01*
X-0014974Y-0023915D02*
Y-0027261D01*
X-0015008Y-0023963D02*
Y-0027261D01*
X-0015043Y-0024010D02*
Y-0027261D01*
X-0015078Y-0024057D02*
Y-0027261D01*
X-0015112Y-0024105D02*
Y-0027261D01*
X-0015147Y-0024152D02*
Y-0027261D01*
X-0015182Y-0024200D02*
Y-0027261D01*
X-0015217Y-0024247D02*
Y-0027261D01*
X-0015251Y-0024294D02*
Y-0027261D01*
X-0015286Y-0024342D02*
Y-0027261D01*
X-0015320Y-0024389D02*
Y-0027261D01*
X-0015355Y-0024437D02*
Y-0027261D01*
X-0015390Y-0024484D02*
Y-0027261D01*
X-0015425Y-0024531D02*
Y-0027261D01*
X-0015459Y-0024579D02*
Y-0027261D01*
X-0015494Y-0024626D02*
Y-0027261D01*
X-0015529Y-0024674D02*
Y-0027261D01*
X-0015563Y-0024721D02*
Y-0027261D01*
X-0015598Y-0024769D02*
Y-0027261D01*
X-0015633Y-0024816D02*
Y-0027261D01*
X-0015667Y-0024863D02*
Y-0027261D01*
X-0015702Y-0024911D02*
Y-0027261D01*
X-0015737Y-0024958D02*
Y-0027261D01*
X-0015772Y-0025006D02*
Y-0027261D01*
X-0015806Y-0025053D02*
Y-0027261D01*
X-0015841Y-0025100D02*
Y-0027261D01*
X-0015876Y-0025148D02*
Y-0027261D01*
X-0015910Y-0025195D02*
Y-0027261D01*
X-0015945Y-0025243D02*
Y-0027261D01*
X-0015980Y-0025290D02*
Y-0027261D01*
X-0016015Y-0025337D02*
Y-0027261D01*
X-0016049Y-0025385D02*
Y-0027261D01*
X-0016084Y-0025432D02*
Y-0027261D01*
X-0016119Y-0025480D02*
Y-0027261D01*
X-0016153Y-0025527D02*
Y-0027261D01*
X-0016188Y-0025574D02*
Y-0027261D01*
X-0016222Y-0025622D02*
Y-0027261D01*
X-0016257Y-0025669D02*
Y-0027261D01*
X-0016292Y-0025717D02*
Y-0027261D01*
X-0016327Y-0025764D02*
Y-0027261D01*
X-0016361Y-0025811D02*
Y-0027261D01*
X-0016396Y-0025859D02*
Y-0027261D01*
X-0016431Y-0025906D02*
Y-0027261D01*
X-0016465Y-0025954D02*
Y-0027261D01*
X-0016500Y-0026001D02*
Y-0027261D01*
X-0016535Y-0026048D02*
Y-0027261D01*
X-0016570Y-0026096D02*
Y-0027261D01*
X-0016604Y-0026143D02*
Y-0027261D01*
X-0016639Y-0026191D02*
Y-0027261D01*
X-0016674Y-0026238D02*
Y-0027261D01*
X-0016708Y-0026285D02*
Y-0027261D01*
X-0016743Y-0026333D02*
Y-0027261D01*
X-0016778Y-0026380D02*
Y-0027261D01*
X-0016813Y-0026428D02*
Y-0027261D01*
X-0016847Y-0026475D02*
Y-0027261D01*
X-0016882Y-0026522D02*
Y-0027261D01*
X-0016917Y-0026570D02*
Y-0027261D01*
X-0016951Y-0026617D02*
Y-0027261D01*
X-0016986Y-0026665D02*
Y-0027261D01*
X-0017020Y-0026712D02*
Y-0027261D01*
X-0017055Y-0026759D02*
Y-0027261D01*
X-0017090Y-0026807D02*
Y-0027261D01*
X-0017125Y-0026854D02*
Y-0027261D01*
X-0017159Y-0026902D02*
Y-0027261D01*
X-0017194Y-0026949D02*
Y-0027261D01*
X-0017229Y-0026996D02*
Y-0027261D01*
X-0017263Y-0027044D02*
Y-0027261D01*
X-0017298Y-0027091D02*
Y-0027261D01*
X-0017333Y-0027139D02*
Y-0027261D01*
X-0017368Y-0027186D02*
Y-0027261D01*
X-0017402Y-0027233D02*
Y-0027261D01*
X-0014252Y-0019192D02*
X-0016834D01*
X-0014232Y-0019226D02*
X-0016811D01*
X-0014211Y-0019261D02*
X-0016787D01*
X-0014191Y-0019296D02*
X-0016763D01*
X-0014170Y-0019330D02*
X-0016739D01*
X-0014150Y-0019365D02*
X-0016715D01*
X-0014130Y-0019400D02*
X-0016691D01*
X-0014109Y-0019435D02*
X-0016668D01*
X-0014089Y-0019469D02*
X-0016644D01*
X-0014068Y-0019504D02*
X-0016620D01*
X-0014048Y-0019539D02*
X-0016596D01*
X-0014027Y-0019573D02*
X-0016572D01*
X-0014007Y-0019608D02*
X-0016548D01*
X-0013986Y-0019643D02*
X-0016525D01*
X-0013966Y-0019677D02*
X-0016501D01*
X-0013945Y-0019712D02*
X-0016477D01*
X-0013925Y-0019747D02*
X-0016453D01*
X-0013904Y-0019781D02*
X-0016430D01*
X-0013884Y-0019816D02*
X-0016406D01*
X-0013864Y-0019851D02*
X-0016382D01*
X-0013843Y-0019885D02*
X-0016358D01*
X-0013823Y-0019920D02*
X-0016334D01*
X-0013802Y-0019955D02*
X-0016310D01*
X-0013782Y-0019990D02*
X-0016287D01*
X-0013761Y-0020024D02*
X-0016263D01*
X-0013741Y-0020059D02*
X-0016239D01*
X-0013720Y-0020094D02*
X-0016215D01*
X-0013700Y-0020128D02*
X-0016191D01*
X-0013680Y-0020163D02*
X-0016167D01*
X-0013659Y-0020198D02*
X-0016144D01*
X-0013639Y-0020232D02*
X-0016120D01*
X-0013618Y-0020267D02*
X-0016096D01*
X-0013598Y-0020302D02*
X-0016072D01*
X-0013577Y-0020337D02*
X-0016048D01*
X-0013557Y-0020371D02*
X-0016024D01*
X-0013536Y-0020406D02*
X-0016001D01*
X-0013516Y-0020441D02*
X-0015977D01*
X-0013495Y-0020475D02*
X-0015953D01*
X-0013475Y-0020510D02*
X-0015929D01*
X-0013454Y-0020545D02*
X-0015906D01*
X-0013434Y-0020580D02*
X-0015881D01*
X-0013413Y-0020614D02*
X-0015858D01*
X-0013393Y-0020649D02*
X-0015834D01*
X-0013373Y-0020683D02*
X-0015810D01*
X-0013352Y-0020718D02*
X-0015786D01*
X-0013332Y-0020753D02*
X-0015763D01*
X-0013311Y-0020787D02*
X-0015739D01*
X-0013291Y-0020822D02*
X-0015715D01*
X-0013270Y-0020857D02*
X-0015691D01*
X-0013250Y-0020892D02*
X-0015667D01*
X-0013230Y-0020926D02*
X-0015643D01*
X-0013209Y-0020961D02*
X-0015620D01*
X-0013189Y-0020996D02*
X-0015596D01*
X-0013168Y-0021030D02*
X-0015572D01*
X-0013148Y-0021065D02*
X-0015548D01*
X-0013127Y-0021100D02*
X-0015524D01*
X-0013107Y-0021135D02*
X-0015500D01*
X-0013086Y-0021169D02*
X-0015477D01*
X-0013066Y-0021204D02*
X-0015453D01*
X-0013045Y-0021239D02*
X-0015429D01*
X-0010650Y-0021273D02*
X-0015405D01*
X-0010674Y-0021308D02*
X-0015381D01*
X-0010698Y-0021343D02*
X-0015357D01*
X-0010721Y-0021378D02*
X-0015334D01*
X-0010745Y-0021412D02*
X-0015310D01*
X-0010769Y-0021447D02*
X-0015286D01*
X-0010793Y-0021481D02*
X-0015262D01*
X-0010817Y-0021516D02*
X-0015239D01*
X-0010841Y-0021551D02*
X-0015215D01*
X-0010865Y-0021585D02*
X-0015191D01*
X-0010888Y-0021620D02*
X-0015167D01*
X-0010912Y-0021655D02*
X-0015143D01*
X-0010936Y-0021690D02*
X-0015119D01*
X-0010960Y-0021724D02*
X-0015096D01*
X-0010983Y-0021759D02*
X-0015072D01*
X-0011007Y-0021794D02*
X-0015048D01*
X-0011031Y-0021828D02*
X-0015024D01*
X-0011055Y-0021863D02*
X-0015000D01*
X-0011079Y-0021898D02*
X-0014976D01*
X-0011103Y-0021933D02*
X-0014953D01*
X-0011126Y-0021967D02*
X-0014929D01*
X-0011150Y-0022002D02*
X-0014905D01*
X-0011174Y-0022037D02*
X-0014881D01*
X-0011198Y-0022071D02*
X-0014857D01*
X-0011222Y-0022106D02*
X-0014833D01*
X-0011246Y-0022141D02*
X-0014810D01*
X-0011269Y-0022175D02*
X-0014786D01*
X-0011293Y-0022210D02*
X-0014762D01*
X-0011317Y-0022245D02*
X-0014738D01*
X-0011341Y-0022280D02*
X-0014715D01*
X-0011365Y-0022314D02*
X-0014691D01*
X-0011389Y-0022349D02*
X-0014667D01*
X-0011412Y-0022383D02*
X-0014643D01*
X-0011436Y-0022418D02*
X-0014619D01*
X-0011460Y-0022453D02*
X-0014595D01*
X-0011484Y-0022488D02*
X-0014572D01*
X-0011508Y-0022522D02*
X-0014548D01*
X-0011531Y-0022557D02*
X-0014524D01*
X-0011556Y-0022592D02*
X-0014500D01*
X-0011579Y-0022626D02*
X-0014476D01*
X-0011603Y-0022661D02*
X-0014452D01*
X-0011627Y-0022696D02*
X-0014429D01*
X-0011651Y-0022730D02*
X-0014405D01*
X-0011674Y-0022765D02*
X-0014381D01*
X-0011698Y-0022800D02*
X-0014357D01*
X-0011722Y-0022835D02*
X-0014333D01*
X-0011746Y-0022869D02*
X-0014309D01*
X-0011770Y-0022904D02*
X-0014286D01*
X-0011794Y-0022939D02*
X-0014262D01*
X-0011772Y-0022973D02*
X-0014284D01*
X-0011748Y-0023008D02*
X-0014310D01*
X-0011724Y-0023043D02*
X-0014335D01*
X-0011700Y-0023078D02*
X-0014361D01*
X-0011676Y-0023112D02*
X-0014386D01*
X-0011652Y-0023147D02*
X-0014411D01*
X-0011628Y-0023181D02*
X-0014437D01*
X-0011604Y-0023216D02*
X-0014462D01*
X-0011580Y-0023251D02*
X-0014487D01*
X-0011556Y-0023285D02*
X-0014513D01*
X-0011532Y-0023320D02*
X-0014538D01*
X-0011508Y-0023355D02*
X-0014564D01*
X-0011484Y-0023390D02*
X-0014589D01*
X-0011460Y-0023424D02*
X-0014615D01*
X-0011436Y-0023459D02*
X-0014640D01*
X-0011412Y-0023494D02*
X-0014665D01*
X-0011388Y-0023528D02*
X-0014691D01*
X-0011364Y-0023563D02*
X-0014716D01*
X-0011340Y-0023598D02*
X-0014741D01*
X-0011316Y-0023633D02*
X-0014767D01*
X-0011292Y-0023667D02*
X-0014792D01*
X-0011268Y-0023702D02*
X-0014818D01*
X-0011244Y-0023737D02*
X-0014843D01*
X-0011220Y-0023771D02*
X-0014869D01*
X-0011196Y-0023806D02*
X-0014894D01*
X-0011172Y-0023841D02*
X-0014919D01*
X-0011148Y-0023876D02*
X-0014944D01*
X-0011124Y-0023910D02*
X-0014970D01*
X-0011100Y-0023945D02*
X-0014995D01*
X-0011076Y-0023980D02*
X-0015021D01*
X-0011052Y-0024014D02*
X-0015046D01*
X-0011028Y-0024049D02*
X-0015072D01*
X-0011004Y-0024083D02*
X-0015097D01*
X-0010980Y-0024118D02*
X-0015122D01*
X-0010956Y-0024153D02*
X-0015148D01*
X-0010932Y-0024188D02*
X-0015173D01*
X-0010908Y-0024222D02*
X-0015198D01*
X-0010884Y-0024257D02*
X-0015224D01*
X-0010860Y-0024292D02*
X-0015249D01*
X-0010836Y-0024326D02*
X-0015275D01*
X-0010812Y-0024361D02*
X-0015300D01*
X-0010788Y-0024396D02*
X-0015326D01*
X-0010764Y-0024431D02*
X-0015351D01*
X-0010740Y-0024465D02*
X-0015376D01*
X-0010716Y-0024500D02*
X-0015402D01*
X-0010692Y-0024535D02*
X-0015427D01*
X-0010668Y-0024569D02*
X-0015452D01*
X-0010644Y-0024604D02*
X-0015478D01*
X-0013037Y-0024639D02*
X-0015503D01*
X-0013062Y-0024673D02*
X-0015529D01*
X-0013086Y-0024708D02*
X-0015554D01*
X-0013111Y-0024743D02*
X-0015580D01*
X-0013135Y-0024778D02*
X-0015605D01*
X-0013159Y-0024812D02*
X-0015630D01*
X-0013184Y-0024847D02*
X-0015656D01*
X-0013208Y-0024881D02*
X-0015681D01*
X-0013233Y-0024916D02*
X-0015706D01*
X-0013257Y-0024951D02*
X-0015732D01*
X-0013281Y-0024986D02*
X-0015757D01*
X-0013306Y-0025020D02*
X-0015783D01*
X-0013330Y-0025055D02*
X-0015808D01*
X-0013355Y-0025090D02*
X-0015833D01*
X-0013379Y-0025124D02*
X-0015859D01*
X-0013404Y-0025159D02*
X-0015884D01*
X-0013428Y-0025194D02*
X-0015909D01*
X-0013452Y-0025228D02*
X-0015935D01*
X-0013477Y-0025263D02*
X-0015960D01*
X-0013501Y-0025298D02*
X-0015986D01*
X-0013526Y-0025333D02*
X-0016011D01*
X-0013550Y-0025367D02*
X-0016037D01*
X-0013574Y-0025402D02*
X-0016062D01*
X-0013599Y-0025437D02*
X-0016087D01*
X-0013623Y-0025471D02*
X-0016113D01*
X-0013648Y-0025506D02*
X-0016138D01*
X-0013672Y-0025541D02*
X-0016163D01*
X-0013696Y-0025576D02*
X-0016189D01*
X-0013721Y-0025610D02*
X-0016214D01*
X-0013745Y-0025645D02*
X-0016240D01*
X-0013770Y-0025680D02*
X-0016265D01*
X-0013794Y-0025714D02*
X-0016291D01*
X-0013819Y-0025749D02*
X-0016316D01*
X-0013843Y-0025783D02*
X-0016341D01*
X-0013867Y-0025819D02*
X-0016367D01*
X-0013892Y-0025853D02*
X-0016392D01*
X-0013916Y-0025888D02*
X-0016417D01*
X-0013941Y-0025922D02*
X-0016443D01*
X-0013965Y-0025957D02*
X-0016468D01*
X-0013989Y-0025992D02*
X-0016494D01*
X-0014014Y-0026026D02*
X-0016519D01*
X-0014038Y-0026061D02*
X-0016544D01*
X-0014063Y-0026096D02*
X-0016570D01*
X-0014087Y-0026131D02*
X-0016595D01*
X-0014111Y-0026165D02*
X-0016620D01*
X-0014136Y-0026200D02*
X-0016646D01*
X-0014160Y-0026235D02*
X-0016671D01*
X-0014185Y-0026269D02*
X-0016697D01*
X-0014209Y-0026304D02*
X-0016722D01*
X-0014233Y-0026339D02*
X-0016748D01*
X-0014258Y-0026374D02*
X-0016773D01*
X-0014282Y-0026408D02*
X-0016798D01*
X-0014307Y-0026443D02*
X-0016824D01*
X-0014331Y-0026478D02*
X-0016849D01*
X-0014356Y-0026512D02*
X-0016874D01*
X-0014380Y-0026547D02*
X-0016900D01*
X-0014404Y-0026581D02*
X-0016925D01*
X-0014429Y-0026616D02*
X-0016951D01*
X-0014453Y-0026651D02*
X-0016976D01*
X-0014478Y-0026686D02*
X-0017002D01*
X-0014502Y-0026720D02*
X-0017027D01*
X-0014526Y-0026755D02*
X-0017052D01*
X-0014551Y-0026790D02*
X-0017078D01*
X-0014575Y-0026824D02*
X-0017103D01*
X-0014600Y-0026859D02*
X-0017128D01*
X-0014624Y-0026894D02*
X-0017154D01*
X-0014648Y-0026929D02*
X-0017179D01*
X-0014673Y-0026963D02*
X-0017205D01*
X-0014697Y-0026998D02*
X-0017230D01*
X-0014722Y-0027033D02*
X-0017256D01*
X-0014746Y-0027067D02*
X-0017281D01*
X-0014770Y-0027102D02*
X-0017306D01*
X-0014795Y-0027137D02*
X-0017331D01*
X-0014819Y-0027171D02*
X-0017357D01*
X-0014844Y-0027206D02*
X-0017382D01*
X-0009249Y-0019178D02*
Y-0019233D01*
X-0009283Y-0019178D02*
Y-0019284D01*
X-0009319Y-0019178D02*
Y-0019334D01*
X-0009353Y-0019178D02*
Y-0019385D01*
X-0009388Y-0019178D02*
Y-0019435D01*
X-0009422Y-0019178D02*
Y-0019486D01*
X-0009457Y-0019178D02*
Y-0019536D01*
X-0009492Y-0019178D02*
Y-0019587D01*
X-0009526Y-0019178D02*
Y-0019637D01*
X-0009561Y-0019178D02*
Y-0019688D01*
X-0009596Y-0019178D02*
Y-0019739D01*
X-0009631Y-0019178D02*
Y-0019789D01*
X-0009665Y-0019178D02*
Y-0019839D01*
X-0009700Y-0019178D02*
Y-0019890D01*
X-0009735Y-0019178D02*
Y-0019941D01*
X-0009769Y-0019178D02*
Y-0019991D01*
X-0009804Y-0019178D02*
Y-0020042D01*
X-0009839Y-0019178D02*
Y-0020092D01*
X-0009874Y-0019178D02*
Y-0020143D01*
X-0009908Y-0019178D02*
Y-0020193D01*
X-0009943Y-0019178D02*
Y-0020244D01*
X-0009978Y-0019178D02*
Y-0020294D01*
X-0010012Y-0019178D02*
Y-0020344D01*
X-0010047Y-0019178D02*
Y-0020395D01*
X-0010081Y-0019178D02*
Y-0020446D01*
X-0010116Y-0019178D02*
Y-0020496D01*
X-0010151Y-0019178D02*
Y-0020547D01*
X-0010186Y-0019178D02*
Y-0020597D01*
X-0010220Y-0019178D02*
Y-0020648D01*
X-0010255Y-0019178D02*
Y-0020698D01*
X-0010290Y-0019178D02*
Y-0020749D01*
X-0010324Y-0019178D02*
Y-0020799D01*
X-0010359Y-0019178D02*
Y-0020850D01*
X-0010394Y-0019178D02*
Y-0020900D01*
X-0010429Y-0019178D02*
Y-0020951D01*
G54D159*
G01X-0009837Y-0034730D02*
X-0010034Y-0034926D01*
Y-0034533D01*
X-0009837Y-0034730D01*
G54D160*
G01X0036474Y-0033086D02*
X0035466D01*
X0035970D02*
Y-0030061D01*
X0035466Y-0030565D01*
X0032944Y-0033086D02*
X0032693Y-0032582D01*
Y-0030565D01*
X0032944Y-0030061D01*
X0034457D01*
X0034709Y-0030565D01*
Y-0032582D01*
X0034457Y-0033086D01*
X0032944D01*
X0031431Y-0031574D02*
X0032440D01*
Y-0032582D01*
X0032187Y-0033086D01*
X0030675D01*
X0030423Y-0032582D01*
Y-0030565D01*
X0030675Y-0030061D01*
X0032187D01*
X0032440Y-0030565D01*
X0028406Y-0033086D02*
X0028154Y-0032582D01*
Y-0030565D01*
X0028406Y-0030061D01*
X0029918D01*
X0030170Y-0030565D01*
Y-0032582D01*
X0029918Y-0033086D01*
X0028406D01*
X0027901D02*
X0026137D01*
Y-0030061D01*
G54D10*
X-0022756Y-0024449D03*
Y-0021220D03*
X-0017913Y-0027854D03*
X-0018386Y-0025886D03*
X-0007559Y-0032047D03*
X-0009528D03*
G54D11*
X-0006575Y-0025591D03*
X-0010512D03*
G54D12*
X0022047Y0028425D03*
X0021260D03*
X-0021260D03*
X-0022047D03*
G54D13*
X0016614Y-0030630D03*
X0016594Y-0031665D03*
Y-0032665D03*
Y-0033665D03*
Y-0034665D03*
X-0020252Y-0019567D03*
X-0019252D03*
X-0018252D03*
X-0022252D03*
X0006508Y-0018059D03*
Y-0019059D03*
Y-0020059D03*
Y-0021059D03*
Y-0022059D03*
Y-0023059D03*
X-0023126Y0026760D03*
X-0022126Y0025760D03*
X-0023126D03*
X-0022126Y0024760D03*
X-0023126D03*
X-0022126Y0023760D03*
X-0023126D03*
X-0022126Y0022760D03*
X-0023126D03*
X-0022126Y0021760D03*
X-0023126D03*
X-0022126Y0020760D03*
X-0023126D03*
X-0022126Y0019760D03*
X-0023126D03*
X-0022126Y0018760D03*
X-0023126D03*
X-0022126Y0017760D03*
X-0023126D03*
X-0022126Y0016760D03*
X-0023126D03*
X-0022126Y0015760D03*
X-0023126D03*
X-0022126Y0014760D03*
X-0023126D03*
X-0022126Y0013760D03*
X-0023126D03*
X-0022126Y0012760D03*
X-0023126D03*
X-0022126Y0011760D03*
X-0023126D03*
X-0022126Y0010760D03*
X-0023126D03*
X-0022126Y0009760D03*
X-0023126D03*
X-0022126Y0008760D03*
X-0023126D03*
X-0022126Y0007760D03*
X-0023126D03*
X-0022126Y0006760D03*
X-0023126D03*
X-0022126Y0005760D03*
X-0023126D03*
X-0022126Y0004760D03*
X-0023126D03*
X-0022126Y0003760D03*
X-0023126D03*
X-0022126Y0002760D03*
X-0023126D03*
X-0022126Y0001768D03*
X-0023126Y0001760D03*
X-0022126Y0000760D03*
X-0023126D03*
X-0022126Y-0000240D03*
X-0023126D03*
X-0022126Y-0001240D03*
X-0023126D03*
X-0022126Y-0002240D03*
X-0023126D03*
X-0022126Y-0003240D03*
X-0023126D03*
X-0022126Y-0004240D03*
X-0023126D03*
X0023126D03*
X0022126Y-0003240D03*
X0023126D03*
X0022126Y-0002240D03*
X0023126D03*
X0022126Y-0001240D03*
X0023126D03*
X0022126Y-0000240D03*
X0023126D03*
X0022126Y0000760D03*
X0023126D03*
X0022126Y0001760D03*
X0023126D03*
X0022126Y0002760D03*
X0023126D03*
X0022126Y0003760D03*
X0023126D03*
X0022126Y0004760D03*
X0023126D03*
X0022126Y0005760D03*
X0023126D03*
X0022126Y0006760D03*
X0023126D03*
X0022126Y0007760D03*
X0023126D03*
X0022126Y0008760D03*
X0023126D03*
X0022126Y0009760D03*
X0023126D03*
X0022126Y0010760D03*
X0023126D03*
X0022126Y0011760D03*
X0023126D03*
X0022126Y0012760D03*
X0023126D03*
X0022126Y0013760D03*
X0023126D03*
X0022126Y0014760D03*
X0023126D03*
X0022126Y0015760D03*
X0023126D03*
X0022126Y0016760D03*
X0023126D03*
X0022126Y0017760D03*
X0023126D03*
X0022126Y0018760D03*
X0023126D03*
X0022126Y0019760D03*
X0023126D03*
X0022126Y0020752D03*
X0023126Y0020760D03*
X0022126Y0021760D03*
X0023126D03*
X0022126Y0022760D03*
X0023126D03*
X0022126Y0023760D03*
X0023126D03*
X0022126Y0024760D03*
X0023126D03*
X0022126Y0025760D03*
X0023126D03*
X0022126Y0026760D03*
X0023126D03*
X0007933Y-0020705D03*
Y-0021705D03*
X-0008063Y-0034717D03*
X-0000969Y0028031D03*
X0000031D03*
X0001031D03*
X0002041D03*
G54D14*
X0016594Y-0029665D03*
X0006508Y-0017059D03*
X-0022126Y0026760D03*
X0022126Y-0004240D03*
X0007933Y-0019705D03*
X-0009063Y-0034717D03*
X-0001969Y0028031D03*
G54D15*
X-0022756Y-0023622D03*
Y-0022835D03*
Y-0022047D03*
X-0005581Y0029846D03*
X-0006081Y0030846D03*
X-0005081D03*
X-0004081D03*
X-0004581Y0029846D03*
X-0003581D03*
X-0002581D03*
X-0003081Y0030846D03*
X-0006941Y0034945D03*
X-0005941D03*
X-0002720D03*
X-0001720D03*
X0003081Y0029846D03*
X0002581Y0030846D03*
X0003581D03*
X0004581D03*
X0004081Y0029846D03*
X0005081D03*
X0006081D03*
X0005581Y0030846D03*
X0001720Y0034945D03*
X0002720D03*
X0005941D03*
X0006941D03*
G54D16*
X-0001281Y0032146D03*
X-0007380D03*
X0007380D03*
X0001281D03*
G54D17*
X-0002081Y0033346D03*
X-0006581D03*
X0006581D03*
X0002081D03*
G54D18*
X0015611Y0027047D03*
X0016319D03*
X0017696D03*
X0016989D03*
X-0006594Y0004843D03*
X-0005886D03*
X-0004508D03*
X-0005216D03*
X-0017696D03*
X-0016989D03*
X-0015611D03*
X-0016319D03*
X0004508D03*
X0005216D03*
X0006594D03*
X0005886D03*
X0015611D03*
X0016319D03*
X0017696D03*
X0016989D03*
X-0006594Y-0006260D03*
X-0005886D03*
X-0004508D03*
X-0005216D03*
X-0017696D03*
X-0016989D03*
X-0015611D03*
X-0016319D03*
X0004508D03*
X0005216D03*
X0006594D03*
X0005886D03*
X0015611D03*
X0016319D03*
X0017696D03*
X0016989D03*
X-0006594Y0015945D03*
X-0005886D03*
X-0004508D03*
X-0005216D03*
X-0017696D03*
X-0016989D03*
X-0015611D03*
X-0016319D03*
X0004508D03*
X0005216D03*
X0006594D03*
X0005886D03*
X0015611D03*
X0016319D03*
X0017696D03*
X0016989D03*
X-0006594Y0027047D03*
X-0005886D03*
X-0004508D03*
X-0005216D03*
X-0017696D03*
X-0016989D03*
X-0015611D03*
X-0016319D03*
X0004508D03*
X0005216D03*
X0006594D03*
X0005886D03*
G54D19*
X0019047Y-0030858D03*
X-0019047D03*
X0019047Y0030858D03*
X-0019047D03*
G54D20*
X-0020571Y-0025118D03*
G54D21*
X-0021752Y-0026969D03*
G54D22*
X-0019390D03*
G54D25*
X-0009173Y0003720D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0003406D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0003091D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0002776D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0002461D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0002146D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0001831D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0001516D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0001201D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0000886D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0000571D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0000256D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0000059D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0000374D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0000689D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0001004D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0001319D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0001634D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0001949D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0002264D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0002579D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0002894D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0003209D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0003524D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0020276Y0003720D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0003406D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0003091D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0002776D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0002461D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0002146D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0001831D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0001516D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0001201D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0000886D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0000571D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0000256D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0000059D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0000374D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0000689D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0001004D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0001319D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0001634D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0001949D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0002264D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0002579D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0002894D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0003209D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0003524D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X0001929Y0003720D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0003406D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0003091D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0002776D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0002461D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0002146D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0001831D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0001516D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0001201D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0000886D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0000571D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0000256D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0000059D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0000374D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0000689D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0001004D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0001319D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0001634D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0001949D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0002264D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0002579D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0002894D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0003209D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0003524D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0013031Y0003720D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0003406D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0003091D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0002776D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0002461D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0002146D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0001831D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0001516D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0001201D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0000886D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0000571D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0000256D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0000059D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0000374D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0000689D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0001004D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0001319D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0001634D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0001949D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0002264D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0002579D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0002894D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0003209D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0003524D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X-0009173Y-0007382D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0007697D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0008012D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0008327D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0008642D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0008957D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0009272D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0009587D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0009902D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0010217D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0010531D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0010846D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0011161D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0011476D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0011791D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0012106D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0012421D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0012736D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0013051D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0013366D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0013681D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0013996D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0014311D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y-0014626D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0020276Y-0007382D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0007697D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0008012D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0008327D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0008642D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0008957D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0009272D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0009587D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0009902D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0010217D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0010531D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0010846D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0011161D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0011476D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0011791D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0012106D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0012421D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0012736D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0013051D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0013366D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0013681D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0013996D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0014311D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y-0014626D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X0001929Y-0007382D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0007697D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0008012D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0008327D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0008642D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0008957D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0009272D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0009587D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0009902D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0010217D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0010531D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0010846D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0011161D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0011476D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0011791D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0012106D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0012421D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0012736D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0013051D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0013366D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0013681D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0013996D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0014311D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y-0014626D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0013031Y-0007382D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0007697D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0008012D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0008327D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0008642D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0008957D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0009272D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0009587D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0009902D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0010217D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0010531D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0010846D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0011161D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0011476D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0011791D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0012106D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0012421D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0012736D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0013051D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0013366D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0013681D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0013996D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0014311D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y-0014626D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X-0009173Y0014823D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0014508D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0014193D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0013878D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0013563D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0013248D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0012933D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0012618D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0012303D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0011988D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0011673D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0011358D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0011043D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0010728D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0010413D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0010098D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0009783D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0009469D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0009154D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0008839D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0008524D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0008209D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0007894D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0007579D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0020276Y0014823D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0014508D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0014193D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0013878D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0013563D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0013248D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0012933D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0012618D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0012303D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0011988D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0011673D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0011358D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0011043D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0010728D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0010413D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0010098D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0009783D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0009469D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0009154D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0008839D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0008524D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0008209D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0007894D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0007579D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X0001929Y0014823D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0014508D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0014193D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0013878D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0013563D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0013248D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0012933D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0012618D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0012303D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0011988D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0011673D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0011358D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0011043D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0010728D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0010413D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0010098D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0009783D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0009469D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0009154D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0008839D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0008524D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0008209D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0007894D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0007579D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0013031Y0014823D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0014508D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0014193D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0013878D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0013563D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0013248D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0012933D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0012618D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0012303D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0011988D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0011673D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0011358D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0011043D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0010728D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0010413D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0010098D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0009783D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0009469D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0009154D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0008839D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0008524D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0008209D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0007894D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0007579D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X-0009173Y0025925D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0025610D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0025295D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0024980D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0024665D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0024350D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0024035D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0023720D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0023406D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0023091D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0022776D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0022461D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0022146D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0021831D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0021516D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0021201D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0020886D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0020571D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0020256D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0019941D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0019626D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0019311D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0018996D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0009173Y0018681D03*
X-0008858D03*
X-0008543D03*
X-0008228D03*
X-0007913D03*
X-0007598D03*
X-0007283D03*
X-0006969D03*
X-0006654D03*
X-0006339D03*
X-0006024D03*
X-0005709D03*
X-0005394D03*
X-0005079D03*
X-0004764D03*
X-0004449D03*
X-0004134D03*
X-0003819D03*
X-0003504D03*
X-0003189D03*
X-0002874D03*
X-0002559D03*
X-0002244D03*
X-0001929D03*
X-0020276Y0025925D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0025610D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0025295D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0024980D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0024665D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0024350D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0024035D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0023720D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0023406D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0023091D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0022776D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0022461D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0022146D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0021831D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0021516D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0021201D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0020886D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0020571D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0020256D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0019941D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0019626D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0019311D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0018996D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X-0020276Y0018681D03*
X-0019961D03*
X-0019646D03*
X-0019331D03*
X-0019016D03*
X-0018701D03*
X-0018386D03*
X-0018071D03*
X-0017756D03*
X-0017441D03*
X-0017126D03*
X-0016811D03*
X-0016496D03*
X-0016181D03*
X-0015866D03*
X-0015551D03*
X-0015236D03*
X-0014921D03*
X-0014606D03*
X-0014291D03*
X-0013976D03*
X-0013661D03*
X-0013346D03*
X-0013031D03*
X0001929Y0025925D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0025610D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0025295D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0024980D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0024665D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0024350D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0024035D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0023720D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0023406D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0023091D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0022776D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0022461D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0022146D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0021831D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0021516D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0021201D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0020886D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0020571D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0020256D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0019941D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0019626D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0019311D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0018996D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0001929Y0018681D03*
X0002244D03*
X0002559D03*
X0002874D03*
X0003189D03*
X0003504D03*
X0003819D03*
X0004134D03*
X0004449D03*
X0004764D03*
X0005079D03*
X0005394D03*
X0005709D03*
X0006024D03*
X0006339D03*
X0006654D03*
X0006969D03*
X0007283D03*
X0007598D03*
X0007913D03*
X0008228D03*
X0008543D03*
X0008858D03*
X0009173D03*
X0013031Y0025925D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0025610D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0025295D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0024980D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0024665D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0024350D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0024035D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0023720D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0023406D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0023091D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0022776D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0022461D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0022146D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0021831D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0021516D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0021201D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0020886D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0020571D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0020256D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0019941D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0019626D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0019311D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0018996D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
X0013031Y0018681D03*
X0013346D03*
X0013661D03*
X0013976D03*
X0014291D03*
X0014606D03*
X0014921D03*
X0015236D03*
X0015551D03*
X0015866D03*
X0016181D03*
X0016496D03*
X0016811D03*
X0017126D03*
X0017441D03*
X0017756D03*
X0018071D03*
X0018386D03*
X0018701D03*
X0019016D03*
X0019331D03*
X0019646D03*
X0019961D03*
X0020276D03*
G54D26*
X-0005453Y-0033307D03*
Y-0029559D03*
Y-0025811D03*
X-0000453Y-0034559D03*
X0000799D03*
X0002051D03*
X0007051D03*
Y-0029559D03*
Y-0028307D03*
Y-0024559D03*
X0002051D03*
X0000799D03*
X-0000453D03*
G54D27*
X0011915Y-0026853D03*
Y-0025603D03*
Y-0024353D03*
X0019415D03*
Y-0028103D03*
G54D28*
X0011915D03*
M02*
